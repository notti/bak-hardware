-------------------------------------------------------------------------------
--$Date: 2008/05/30 00:57:53 $
--$RCSfile: multi_mgt_wrapper_vhd.ejava,v $
--$Revision: 1.1.2.1 $
-------------------------------------------------------------------------------
--   ____  ____ 
--  /   /\/   / 
-- /___/  \  /    Vendor: Xilinx 
-- \   \   \/     Version : 1.5 
--  \   \         Application : RocketIO GTX Wizard 
--  /   /         Filename : gtx.vhd
-- /___/   /\     Timestamp : 02/08/2005 09:12:43
-- \   \  /  \ 
--  \___\/\___\ 
--
--
-- Module GTX (a GTX Wrapper)
-- Generated by Xilinx RocketIO GTX Wizard

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***************************** Entity Declaration ****************************

entity GTX is
generic
(
    -- Simulation attributes
    WRAPPER_SIM_MODE                : string    := "FAST"; -- Set to Fast Functional Simulation Model
    WRAPPER_SIM_GTXRESET_SPEEDUP    : integer   := 0; -- Set to 1 to speed up sim reset
    WRAPPER_SIM_PLL_PERDIV2         : bit_vector:= x"0fa" -- Set to the VCO Unit Interval time
);
port
(
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE0  (Location)

    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    TILE0_RXCHARISCOMMA0_OUT                : out  std_logic_vector(1 downto 0);
    TILE0_RXCHARISCOMMA1_OUT                : out  std_logic_vector(1 downto 0);
    TILE0_RXDISPERR0_OUT                    : out  std_logic_vector(1 downto 0);
    TILE0_RXDISPERR1_OUT                    : out  std_logic_vector(1 downto 0);
    TILE0_RXNOTINTABLE0_OUT                 : out  std_logic_vector(1 downto 0);
    TILE0_RXNOTINTABLE1_OUT                 : out  std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    TILE0_RXBYTEISALIGNED0_OUT              : out  std_logic;
    TILE0_RXBYTEISALIGNED1_OUT              : out  std_logic;
    TILE0_RXBYTEREALIGN0_OUT                : out  std_logic;
    TILE0_RXBYTEREALIGN1_OUT                : out  std_logic;
    TILE0_RXENMCOMMAALIGN0_IN               : in   std_logic;
    TILE0_RXENMCOMMAALIGN1_IN               : in   std_logic;
    TILE0_RXENPCOMMAALIGN0_IN               : in   std_logic;
    TILE0_RXENPCOMMAALIGN1_IN               : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    TILE0_RXDATA0_OUT                       : out  std_logic_vector(15 downto 0);
    TILE0_RXDATA1_OUT                       : out  std_logic_vector(15 downto 0);
    TILE0_RXUSRCLK0_IN                      : in   std_logic;
    TILE0_RXUSRCLK1_IN                      : in   std_logic;
    TILE0_RXUSRCLK20_IN                     : in   std_logic;
    TILE0_RXUSRCLK21_IN                     : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    TILE0_RXEQMIX0_IN                       : in   std_logic_vector(1 downto 0);
    TILE0_RXEQMIX1_IN                       : in   std_logic_vector(1 downto 0);
    TILE0_RXN0_IN                           : in   std_logic;
    TILE0_RXN1_IN                           : in   std_logic;
    TILE0_RXP0_IN                           : in   std_logic;
    TILE0_RXP1_IN                           : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    TILE0_RXPOLARITY0_IN                    : in   std_logic;
    TILE0_RXPOLARITY1_IN                    : in   std_logic;
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    TILE0_CLKIN_IN                          : in   std_logic;
    TILE0_GTXRESET_IN                       : in   std_logic;
    TILE0_PLLLKDET_OUT                      : out  std_logic;
    TILE0_REFCLKOUT_OUT                     : out  std_logic;
    TILE0_RESETDONE0_OUT                    : out  std_logic;
    TILE0_RESETDONE1_OUT                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TILE0_TXDATA0_IN                        : in   std_logic_vector(19 downto 0);
    TILE0_TXDATA1_IN                        : in   std_logic_vector(19 downto 0);
    TILE0_TXUSRCLK0_IN                      : in   std_logic;
    TILE0_TXUSRCLK1_IN                      : in   std_logic;
    TILE0_TXUSRCLK20_IN                     : in   std_logic;
    TILE0_TXUSRCLK21_IN                     : in   std_logic;
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    TILE0_TXN0_OUT                          : out  std_logic;
    TILE0_TXN1_OUT                          : out  std_logic;
    TILE0_TXP0_OUT                          : out  std_logic;
    TILE0_TXP1_OUT                          : out  std_logic;


    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE1  (Location)

    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    TILE1_RXCHARISCOMMA0_OUT                : out  std_logic_vector(1 downto 0);
    TILE1_RXCHARISCOMMA1_OUT                : out  std_logic_vector(1 downto 0);
    TILE1_RXDISPERR0_OUT                    : out  std_logic_vector(1 downto 0);
    TILE1_RXDISPERR1_OUT                    : out  std_logic_vector(1 downto 0);
    TILE1_RXNOTINTABLE0_OUT                 : out  std_logic_vector(1 downto 0);
    TILE1_RXNOTINTABLE1_OUT                 : out  std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    TILE1_RXBYTEISALIGNED0_OUT              : out  std_logic;
    TILE1_RXBYTEISALIGNED1_OUT              : out  std_logic;
    TILE1_RXBYTEREALIGN0_OUT                : out  std_logic;
    TILE1_RXBYTEREALIGN1_OUT                : out  std_logic;
    TILE1_RXENMCOMMAALIGN0_IN               : in   std_logic;
    TILE1_RXENMCOMMAALIGN1_IN               : in   std_logic;
    TILE1_RXENPCOMMAALIGN0_IN               : in   std_logic;
    TILE1_RXENPCOMMAALIGN1_IN               : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    TILE1_RXDATA0_OUT                       : out  std_logic_vector(15 downto 0);
    TILE1_RXDATA1_OUT                       : out  std_logic_vector(15 downto 0);
    TILE1_RXUSRCLK0_IN                      : in   std_logic;
    TILE1_RXUSRCLK1_IN                      : in   std_logic;
    TILE1_RXUSRCLK20_IN                     : in   std_logic;
    TILE1_RXUSRCLK21_IN                     : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    TILE1_RXEQMIX0_IN                       : in   std_logic_vector(1 downto 0);
    TILE1_RXEQMIX1_IN                       : in   std_logic_vector(1 downto 0);
    TILE1_RXN0_IN                           : in   std_logic;
    TILE1_RXN1_IN                           : in   std_logic;
    TILE1_RXP0_IN                           : in   std_logic;
    TILE1_RXP1_IN                           : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    TILE1_RXPOLARITY0_IN                    : in   std_logic;
    TILE1_RXPOLARITY1_IN                    : in   std_logic;
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    TILE1_CLKIN_IN                          : in   std_logic;
    TILE1_GTXRESET_IN                       : in   std_logic;
    TILE1_PLLLKDET_OUT                      : out  std_logic;
    TILE1_REFCLKOUT_OUT                     : out  std_logic;
    TILE1_RESETDONE0_OUT                    : out  std_logic;
    TILE1_RESETDONE1_OUT                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TILE1_TXDATA0_IN                        : in   std_logic_vector(19 downto 0);
    TILE1_TXDATA1_IN                        : in   std_logic_vector(19 downto 0);
    TILE1_TXUSRCLK0_IN                      : in   std_logic;
    TILE1_TXUSRCLK1_IN                      : in   std_logic;
    TILE1_TXUSRCLK20_IN                     : in   std_logic;
    TILE1_TXUSRCLK21_IN                     : in   std_logic;
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    TILE1_TXN0_OUT                          : out  std_logic;
    TILE1_TXN1_OUT                          : out  std_logic;
    TILE1_TXP0_OUT                          : out  std_logic;
    TILE1_TXP1_OUT                          : out  std_logic


);

    attribute X_CORE_INFO : string;
    attribute X_CORE_INFO of GTX : entity is "gtxwizard_v1_5, Coregen v10.1_ip3";

end GTX;

architecture RTL of GTX is

--***************************** Signal Declarations *****************************

    -- Channel Bonding Signals
    signal  tile0_rxchbondo0_i   : std_logic_vector(3 downto 0);
    signal  tile0_rxchbondo1_i   : std_logic_vector(3 downto 0);

    signal  tile1_rxchbondo0_i   : std_logic_vector(3 downto 0);
    signal  tile1_rxchbondo1_i   : std_logic_vector(3 downto 0);


    -- ground and tied_to_vcc_i signals
    signal  tied_to_ground_i                :   std_logic;
    signal  tied_to_ground_vec_i            :   std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   :   std_logic;
    

--*************************** Component Declarations **************************

component GTX_TILE 
generic
(
    -- Simulation attributes
    TILE_SIM_MODE                : string    := "FAST"; -- Set to Fast Functional Simulation Model
    TILE_SIM_GTXRESET_SPEEDUP    : integer   := 0; -- Set to 1 to speed up sim reset
    TILE_SIM_PLL_PERDIV2         : bit_vector:= x"0fa"; -- Set to the VCO Unit Interval time 

    -- Channel bonding attributes
    TILE_CHAN_BOND_MODE_0        : string    := "OFF";  -- "MASTER", "SLAVE", or "OFF"
    TILE_CHAN_BOND_LEVEL_0       : integer   := 0;     -- 0 to 7. See UG for details
    
    TILE_CHAN_BOND_MODE_1        : string    := "OFF";  -- "MASTER", "SLAVE", or "OFF"
    TILE_CHAN_BOND_LEVEL_1       : integer   := 0      -- 0 to 7. See UG for details
);
port 
(   
    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    RXCHARISCOMMA0_OUT                      : out  std_logic_vector(1 downto 0);
    RXCHARISCOMMA1_OUT                      : out  std_logic_vector(1 downto 0);
    RXDISPERR0_OUT                          : out  std_logic_vector(1 downto 0);
    RXDISPERR1_OUT                          : out  std_logic_vector(1 downto 0);
    RXNOTINTABLE0_OUT                       : out  std_logic_vector(1 downto 0);
    RXNOTINTABLE1_OUT                       : out  std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    RXBYTEISALIGNED0_OUT                    : out  std_logic;
    RXBYTEISALIGNED1_OUT                    : out  std_logic;
    RXBYTEREALIGN0_OUT                      : out  std_logic;
    RXBYTEREALIGN1_OUT                      : out  std_logic;
    RXENMCOMMAALIGN0_IN                     : in   std_logic;
    RXENMCOMMAALIGN1_IN                     : in   std_logic;
    RXENPCOMMAALIGN0_IN                     : in   std_logic;
    RXENPCOMMAALIGN1_IN                     : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    RXDATA0_OUT                             : out  std_logic_vector(15 downto 0);
    RXDATA1_OUT                             : out  std_logic_vector(15 downto 0);
    RXUSRCLK0_IN                            : in   std_logic;
    RXUSRCLK1_IN                            : in   std_logic;
    RXUSRCLK20_IN                           : in   std_logic;
    RXUSRCLK21_IN                           : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    RXEQMIX0_IN                             : in   std_logic_vector(1 downto 0);
    RXEQMIX1_IN                             : in   std_logic_vector(1 downto 0);
    RXN0_IN                                 : in   std_logic;
    RXN1_IN                                 : in   std_logic;
    RXP0_IN                                 : in   std_logic;
    RXP1_IN                                 : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    RXPOLARITY0_IN                          : in   std_logic;
    RXPOLARITY1_IN                          : in   std_logic;
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    CLKIN_IN                                : in   std_logic;
    GTXRESET_IN                             : in   std_logic;
    PLLLKDET_OUT                            : out  std_logic;
    REFCLKOUT_OUT                           : out  std_logic;
    RESETDONE0_OUT                          : out  std_logic;
    RESETDONE1_OUT                          : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TXDATA0_IN                              : in   std_logic_vector(19 downto 0);
    TXDATA1_IN                              : in   std_logic_vector(19 downto 0);
    TXUSRCLK0_IN                            : in   std_logic;
    TXUSRCLK1_IN                            : in   std_logic;
    TXUSRCLK20_IN                           : in   std_logic;
    TXUSRCLK21_IN                           : in   std_logic;
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    TXN0_OUT                                : out  std_logic;
    TXN1_OUT                                : out  std_logic;
    TXP0_OUT                                : out  std_logic;
    TXP1_OUT                                : out  std_logic


);
end component;


--********************************* Main Body of Code**************************

begin                       

    tied_to_ground_i                    <= '0';
    tied_to_ground_vec_i(63 downto 0)   <= (others => '0');
    tied_to_vcc_i                       <= '1';

    --------------------------- Tile Instances  -------------------------------   


    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE0  (Location)

    tile0_gtx_i : GTX_TILE
    generic map
    (
        -- Simulation attributes
        TILE_SIM_MODE                => WRAPPER_SIM_MODE,
        TILE_SIM_GTXRESET_SPEEDUP    => WRAPPER_SIM_GTXRESET_SPEEDUP,
        TILE_SIM_PLL_PERDIV2         => WRAPPER_SIM_PLL_PERDIV2,

        -- Channel bonding attributes
        TILE_CHAN_BOND_MODE_0        => "OFF",
        TILE_CHAN_BOND_LEVEL_0       => 0,
    
        TILE_CHAN_BOND_MODE_1        => "OFF",
        TILE_CHAN_BOND_LEVEL_1       => 0
    )
    port map
    (
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISCOMMA0_OUT              =>      TILE0_RXCHARISCOMMA0_OUT,
        RXCHARISCOMMA1_OUT              =>      TILE0_RXCHARISCOMMA1_OUT,
        RXDISPERR0_OUT                  =>      TILE0_RXDISPERR0_OUT,
        RXDISPERR1_OUT                  =>      TILE0_RXDISPERR1_OUT,
        RXNOTINTABLE0_OUT               =>      TILE0_RXNOTINTABLE0_OUT,
        RXNOTINTABLE1_OUT               =>      TILE0_RXNOTINTABLE1_OUT,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED0_OUT            =>      TILE0_RXBYTEISALIGNED0_OUT,
        RXBYTEISALIGNED1_OUT            =>      TILE0_RXBYTEISALIGNED1_OUT,
        RXBYTEREALIGN0_OUT              =>      TILE0_RXBYTEREALIGN0_OUT,
        RXBYTEREALIGN1_OUT              =>      TILE0_RXBYTEREALIGN1_OUT,
        RXENMCOMMAALIGN0_IN             =>      TILE0_RXENMCOMMAALIGN0_IN,
        RXENMCOMMAALIGN1_IN             =>      TILE0_RXENMCOMMAALIGN1_IN,
        RXENPCOMMAALIGN0_IN             =>      TILE0_RXENPCOMMAALIGN0_IN,
        RXENPCOMMAALIGN1_IN             =>      TILE0_RXENPCOMMAALIGN1_IN,
        ------------------- Receive Ports - RX Data Path interface -----------------
        RXDATA0_OUT                     =>      TILE0_RXDATA0_OUT,
        RXDATA1_OUT                     =>      TILE0_RXDATA1_OUT,
        RXUSRCLK0_IN                    =>      TILE0_RXUSRCLK0_IN,
        RXUSRCLK1_IN                    =>      TILE0_RXUSRCLK1_IN,
        RXUSRCLK20_IN                   =>      TILE0_RXUSRCLK20_IN,
        RXUSRCLK21_IN                   =>      TILE0_RXUSRCLK21_IN,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        RXEQMIX0_IN                     =>      TILE0_RXEQMIX0_IN,
        RXEQMIX1_IN                     =>      TILE0_RXEQMIX1_IN,
        RXN0_IN                         =>      TILE0_RXN0_IN,
        RXN1_IN                         =>      TILE0_RXN1_IN,
        RXP0_IN                         =>      TILE0_RXP0_IN,
        RXP1_IN                         =>      TILE0_RXP1_IN,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        RXPOLARITY0_IN                  =>      TILE0_RXPOLARITY0_IN,
        RXPOLARITY1_IN                  =>      TILE0_RXPOLARITY1_IN,
        --------------------- Shared Ports - Tile and PLL Ports --------------------
        CLKIN_IN                        =>      TILE0_CLKIN_IN,
        GTXRESET_IN                     =>      TILE0_GTXRESET_IN,
        PLLLKDET_OUT                    =>      TILE0_PLLLKDET_OUT,
        REFCLKOUT_OUT                   =>      TILE0_REFCLKOUT_OUT,
        RESETDONE0_OUT                  =>      TILE0_RESETDONE0_OUT,
        RESETDONE1_OUT                  =>      TILE0_RESETDONE1_OUT,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA0_IN                      =>      TILE0_TXDATA0_IN,
        TXDATA1_IN                      =>      TILE0_TXDATA1_IN,
        TXUSRCLK0_IN                    =>      TILE0_TXUSRCLK0_IN,
        TXUSRCLK1_IN                    =>      TILE0_TXUSRCLK1_IN,
        TXUSRCLK20_IN                   =>      TILE0_TXUSRCLK20_IN,
        TXUSRCLK21_IN                   =>      TILE0_TXUSRCLK21_IN,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TXN0_OUT                        =>      TILE0_TXN0_OUT,
        TXN1_OUT                        =>      TILE0_TXN1_OUT,
        TXP0_OUT                        =>      TILE0_TXP0_OUT,
        TXP1_OUT                        =>      TILE0_TXP1_OUT

    );


    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE1  (Location)

    tile1_gtx_i : GTX_TILE
    generic map
    (
        -- Simulation attributes
        TILE_SIM_MODE                => WRAPPER_SIM_MODE,
        TILE_SIM_GTXRESET_SPEEDUP    => WRAPPER_SIM_GTXRESET_SPEEDUP,
        TILE_SIM_PLL_PERDIV2         => WRAPPER_SIM_PLL_PERDIV2,

        -- Channel bonding attributes
        TILE_CHAN_BOND_MODE_0        => "OFF",
        TILE_CHAN_BOND_LEVEL_0       => 0,
    
        TILE_CHAN_BOND_MODE_1        => "OFF",
        TILE_CHAN_BOND_LEVEL_1       => 0
    )
    port map
    (
        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        RXCHARISCOMMA0_OUT              =>      TILE1_RXCHARISCOMMA0_OUT,
        RXCHARISCOMMA1_OUT              =>      TILE1_RXCHARISCOMMA1_OUT,
        RXDISPERR0_OUT                  =>      TILE1_RXDISPERR0_OUT,
        RXDISPERR1_OUT                  =>      TILE1_RXDISPERR1_OUT,
        RXNOTINTABLE0_OUT               =>      TILE1_RXNOTINTABLE0_OUT,
        RXNOTINTABLE1_OUT               =>      TILE1_RXNOTINTABLE1_OUT,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        RXBYTEISALIGNED0_OUT            =>      TILE1_RXBYTEISALIGNED0_OUT,
        RXBYTEISALIGNED1_OUT            =>      TILE1_RXBYTEISALIGNED1_OUT,
        RXBYTEREALIGN0_OUT              =>      TILE1_RXBYTEREALIGN0_OUT,
        RXBYTEREALIGN1_OUT              =>      TILE1_RXBYTEREALIGN1_OUT,
        RXENMCOMMAALIGN0_IN             =>      TILE1_RXENMCOMMAALIGN0_IN,
        RXENMCOMMAALIGN1_IN             =>      TILE1_RXENMCOMMAALIGN1_IN,
        RXENPCOMMAALIGN0_IN             =>      TILE1_RXENPCOMMAALIGN0_IN,
        RXENPCOMMAALIGN1_IN             =>      TILE1_RXENPCOMMAALIGN1_IN,
        ------------------- Receive Ports - RX Data Path interface -----------------
        RXDATA0_OUT                     =>      TILE1_RXDATA0_OUT,
        RXDATA1_OUT                     =>      TILE1_RXDATA1_OUT,
        RXUSRCLK0_IN                    =>      TILE1_RXUSRCLK0_IN,
        RXUSRCLK1_IN                    =>      TILE1_RXUSRCLK1_IN,
        RXUSRCLK20_IN                   =>      TILE1_RXUSRCLK20_IN,
        RXUSRCLK21_IN                   =>      TILE1_RXUSRCLK21_IN,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        RXEQMIX0_IN                     =>      TILE1_RXEQMIX0_IN,
        RXEQMIX1_IN                     =>      TILE1_RXEQMIX1_IN,
        RXN0_IN                         =>      TILE1_RXN0_IN,
        RXN1_IN                         =>      TILE1_RXN1_IN,
        RXP0_IN                         =>      TILE1_RXP0_IN,
        RXP1_IN                         =>      TILE1_RXP1_IN,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        RXPOLARITY0_IN                  =>      TILE1_RXPOLARITY0_IN,
        RXPOLARITY1_IN                  =>      TILE1_RXPOLARITY1_IN,
        --------------------- Shared Ports - Tile and PLL Ports --------------------
        CLKIN_IN                        =>      TILE1_CLKIN_IN,
        GTXRESET_IN                     =>      TILE1_GTXRESET_IN,
        PLLLKDET_OUT                    =>      TILE1_PLLLKDET_OUT,
        REFCLKOUT_OUT                   =>      TILE1_REFCLKOUT_OUT,
        RESETDONE0_OUT                  =>      TILE1_RESETDONE0_OUT,
        RESETDONE1_OUT                  =>      TILE1_RESETDONE1_OUT,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TXDATA0_IN                      =>      TILE1_TXDATA0_IN,
        TXDATA1_IN                      =>      TILE1_TXDATA1_IN,
        TXUSRCLK0_IN                    =>      TILE1_TXUSRCLK0_IN,
        TXUSRCLK1_IN                    =>      TILE1_TXUSRCLK1_IN,
        TXUSRCLK20_IN                   =>      TILE1_TXUSRCLK20_IN,
        TXUSRCLK21_IN                   =>      TILE1_TXUSRCLK21_IN,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TXN0_OUT                        =>      TILE1_TXN0_OUT,
        TXN1_OUT                        =>      TILE1_TXN1_OUT,
        TXP0_OUT                        =>      TILE1_TXP0_OUT,
        TXP1_OUT                        =>      TILE1_TXP1_OUT

    );

    
     
end RTL;
