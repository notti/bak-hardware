------------------------------------------------------------------------------
--$Date: 2008/07/23 00:16:39 $
--$RCSfile: example_mgt_top_vhd.ejava,v $
--$Revision: 1.1.2.7 $
------------------------------------------------------------------------------
--   ____  ____ 
--  /   /\/   / 
-- /___/  \  /    Vendor: Xilinx 
-- \   \   \/     Version : 1.5
--  \   \         Application : RocketIO GTX Wizard 
--  /   /         Filename : example_mgt_top.vhd
-- /___/   /\     Timestamp : 
-- \   \  /  \ 
--  \___\/\___\ 
--
--
-- Module EXAMPLE_MGT_TOP
-- Generated by Xilinx RocketIO GTX Wizard

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;



--***********************************Entity Declaration************************

entity EXAMPLE_MGT_TOP is
generic
(
    EXAMPLE_CONFIG_INDEPENDENT_LANES        : integer   := 1;
    EXAMPLE_LANE_WITH_START_CHAR            : integer   := 0;
    EXAMPLE_WORDS_IN_BRAM                   : integer   := 512;
    EXAMPLE_SIM_MODE                        : string    := "FAST";
    EXAMPLE_SIM_GTXRESET_SPEEDUP            : integer   := 1;
    EXAMPLE_SIM_PLL_PERDIV2                 : bit_vector:= x"0fa";
    EXAMPLE_USE_CHIPSCOPE                   : integer   := 1     -- Set to 1 to use Chipscope to drive resets
);
port
(
    TILE2_REFCLK_PAD_N_IN                   : in   std_logic;
    TILE2_REFCLK_PAD_P_IN                   : in   std_logic;
    GTXRESET_IN                             : in   std_logic;
    TILE0_PLLLKDET_OUT                      : out  std_logic;
    TILE1_PLLLKDET_OUT                      : out  std_logic;
    TILE2_PLLLKDET_OUT                      : out  std_logic;
    RXN_IN                                  : in   std_logic_vector(5 downto 0);
    RXP_IN                                  : in   std_logic_vector(5 downto 0);
    TXN_OUT                                 : out  std_logic_vector(5 downto 0);
    TXP_OUT                                 : out  std_logic_vector(5 downto 0)
    
);

    attribute X_CORE_INFO : string;
    attribute X_CORE_INFO of EXAMPLE_MGT_TOP : entity is "gtxwizard_v1_5, Coregen v10.1_ip3";

end EXAMPLE_MGT_TOP;
    
architecture RTL of EXAMPLE_MGT_TOP is

--**************************Component Declarations*****************************


component GTX 
generic
(
    -- Simulation attributes
    WRAPPER_SIM_MODE                : string    := "FAST"; -- Set to Fast Functional Simulation Model
    WRAPPER_SIM_GTXRESET_SPEEDUP    : integer   := 0; -- Set to 1 to speed up sim reset
    WRAPPER_SIM_PLL_PERDIV2         : bit_vector:= x"0fa" -- Set to the VCO Unit Interval time
);
port
(
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE0  (Location)

    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    TILE0_RXCHARISCOMMA0_OUT                : out  std_logic_vector(1 downto 0);
    TILE0_RXCHARISCOMMA1_OUT                : out  std_logic_vector(1 downto 0);
    TILE0_RXDISPERR0_OUT                    : out  std_logic_vector(1 downto 0);
    TILE0_RXDISPERR1_OUT                    : out  std_logic_vector(1 downto 0);
    TILE0_RXNOTINTABLE0_OUT                 : out  std_logic_vector(1 downto 0);
    TILE0_RXNOTINTABLE1_OUT                 : out  std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    TILE0_RXBYTEISALIGNED0_OUT              : out  std_logic;
    TILE0_RXBYTEISALIGNED1_OUT              : out  std_logic;
    TILE0_RXENMCOMMAALIGN0_IN               : in   std_logic;
    TILE0_RXENMCOMMAALIGN1_IN               : in   std_logic;
    TILE0_RXENPCOMMAALIGN0_IN               : in   std_logic;
    TILE0_RXENPCOMMAALIGN1_IN               : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    TILE0_RXDATA0_OUT                       : out  std_logic_vector(15 downto 0);
    TILE0_RXDATA1_OUT                       : out  std_logic_vector(15 downto 0);
    TILE0_RXRECCLK0_OUT                     : out  std_logic;
    TILE0_RXRECCLK1_OUT                     : out  std_logic;
    TILE0_RXUSRCLK0_IN                      : in   std_logic;
    TILE0_RXUSRCLK1_IN                      : in   std_logic;
    TILE0_RXUSRCLK20_IN                     : in   std_logic;
    TILE0_RXUSRCLK21_IN                     : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    TILE0_RXEQMIX0_IN                       : in   std_logic_vector(1 downto 0);
    TILE0_RXEQMIX1_IN                       : in   std_logic_vector(1 downto 0);
    TILE0_RXN0_IN                           : in   std_logic;
    TILE0_RXN1_IN                           : in   std_logic;
    TILE0_RXP0_IN                           : in   std_logic;
    TILE0_RXP1_IN                           : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    TILE0_RXPOLARITY0_IN                    : in   std_logic;
    TILE0_RXPOLARITY1_IN                    : in   std_logic;
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    TILE0_CLKIN_IN                          : in   std_logic;
    TILE0_GTXRESET_IN                       : in   std_logic;
    TILE0_PLLLKDET_OUT                      : out  std_logic;
    TILE0_REFCLKOUT_OUT                     : out  std_logic;
    TILE0_RESETDONE0_OUT                    : out  std_logic;
    TILE0_RESETDONE1_OUT                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TILE0_TXDATA0_IN                        : in   std_logic_vector(19 downto 0);
    TILE0_TXDATA1_IN                        : in   std_logic_vector(19 downto 0);
    TILE0_TXUSRCLK0_IN                      : in   std_logic;
    TILE0_TXUSRCLK1_IN                      : in   std_logic;
    TILE0_TXUSRCLK20_IN                     : in   std_logic;
    TILE0_TXUSRCLK21_IN                     : in   std_logic;
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    TILE0_TXN0_OUT                          : out  std_logic;
    TILE0_TXN1_OUT                          : out  std_logic;
    TILE0_TXP0_OUT                          : out  std_logic;
    TILE0_TXP1_OUT                          : out  std_logic;


    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE1  (Location)

    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    TILE1_RXCHARISCOMMA0_OUT                : out  std_logic_vector(1 downto 0);
    TILE1_RXCHARISCOMMA1_OUT                : out  std_logic_vector(1 downto 0);
    TILE1_RXDISPERR0_OUT                    : out  std_logic_vector(1 downto 0);
    TILE1_RXDISPERR1_OUT                    : out  std_logic_vector(1 downto 0);
    TILE1_RXNOTINTABLE0_OUT                 : out  std_logic_vector(1 downto 0);
    TILE1_RXNOTINTABLE1_OUT                 : out  std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    TILE1_RXBYTEISALIGNED0_OUT              : out  std_logic;
    TILE1_RXBYTEISALIGNED1_OUT              : out  std_logic;
    TILE1_RXENMCOMMAALIGN0_IN               : in   std_logic;
    TILE1_RXENMCOMMAALIGN1_IN               : in   std_logic;
    TILE1_RXENPCOMMAALIGN0_IN               : in   std_logic;
    TILE1_RXENPCOMMAALIGN1_IN               : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    TILE1_RXDATA0_OUT                       : out  std_logic_vector(15 downto 0);
    TILE1_RXDATA1_OUT                       : out  std_logic_vector(15 downto 0);
    TILE1_RXRECCLK0_OUT                     : out  std_logic;
    TILE1_RXRECCLK1_OUT                     : out  std_logic;
    TILE1_RXUSRCLK0_IN                      : in   std_logic;
    TILE1_RXUSRCLK1_IN                      : in   std_logic;
    TILE1_RXUSRCLK20_IN                     : in   std_logic;
    TILE1_RXUSRCLK21_IN                     : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    TILE1_RXEQMIX0_IN                       : in   std_logic_vector(1 downto 0);
    TILE1_RXEQMIX1_IN                       : in   std_logic_vector(1 downto 0);
    TILE1_RXN0_IN                           : in   std_logic;
    TILE1_RXN1_IN                           : in   std_logic;
    TILE1_RXP0_IN                           : in   std_logic;
    TILE1_RXP1_IN                           : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    TILE1_RXPOLARITY0_IN                    : in   std_logic;
    TILE1_RXPOLARITY1_IN                    : in   std_logic;
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    TILE1_CLKIN_IN                          : in   std_logic;
    TILE1_GTXRESET_IN                       : in   std_logic;
    TILE1_PLLLKDET_OUT                      : out  std_logic;
    TILE1_REFCLKOUT_OUT                     : out  std_logic;
    TILE1_RESETDONE0_OUT                    : out  std_logic;
    TILE1_RESETDONE1_OUT                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TILE1_TXDATA0_IN                        : in   std_logic_vector(19 downto 0);
    TILE1_TXDATA1_IN                        : in   std_logic_vector(19 downto 0);
    TILE1_TXUSRCLK0_IN                      : in   std_logic;
    TILE1_TXUSRCLK1_IN                      : in   std_logic;
    TILE1_TXUSRCLK20_IN                     : in   std_logic;
    TILE1_TXUSRCLK21_IN                     : in   std_logic;
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    TILE1_TXN0_OUT                          : out  std_logic;
    TILE1_TXN1_OUT                          : out  std_logic;
    TILE1_TXP0_OUT                          : out  std_logic;
    TILE1_TXP1_OUT                          : out  std_logic;


    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE2  (Location)

    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    TILE2_RXCHARISCOMMA0_OUT                : out  std_logic_vector(1 downto 0);
    TILE2_RXCHARISCOMMA1_OUT                : out  std_logic_vector(1 downto 0);
    TILE2_RXDISPERR0_OUT                    : out  std_logic_vector(1 downto 0);
    TILE2_RXDISPERR1_OUT                    : out  std_logic_vector(1 downto 0);
    TILE2_RXNOTINTABLE0_OUT                 : out  std_logic_vector(1 downto 0);
    TILE2_RXNOTINTABLE1_OUT                 : out  std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    TILE2_RXBYTEISALIGNED0_OUT              : out  std_logic;
    TILE2_RXBYTEISALIGNED1_OUT              : out  std_logic;
    TILE2_RXENMCOMMAALIGN0_IN               : in   std_logic;
    TILE2_RXENMCOMMAALIGN1_IN               : in   std_logic;
    TILE2_RXENPCOMMAALIGN0_IN               : in   std_logic;
    TILE2_RXENPCOMMAALIGN1_IN               : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    TILE2_RXDATA0_OUT                       : out  std_logic_vector(15 downto 0);
    TILE2_RXDATA1_OUT                       : out  std_logic_vector(15 downto 0);
    TILE2_RXRECCLK0_OUT                     : out  std_logic;
    TILE2_RXRECCLK1_OUT                     : out  std_logic;
    TILE2_RXUSRCLK0_IN                      : in   std_logic;
    TILE2_RXUSRCLK1_IN                      : in   std_logic;
    TILE2_RXUSRCLK20_IN                     : in   std_logic;
    TILE2_RXUSRCLK21_IN                     : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    TILE2_RXEQMIX0_IN                       : in   std_logic_vector(1 downto 0);
    TILE2_RXEQMIX1_IN                       : in   std_logic_vector(1 downto 0);
    TILE2_RXN0_IN                           : in   std_logic;
    TILE2_RXN1_IN                           : in   std_logic;
    TILE2_RXP0_IN                           : in   std_logic;
    TILE2_RXP1_IN                           : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    TILE2_RXPOLARITY0_IN                    : in   std_logic;
    TILE2_RXPOLARITY1_IN                    : in   std_logic;
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    TILE2_CLKIN_IN                          : in   std_logic;
    TILE2_GTXRESET_IN                       : in   std_logic;
    TILE2_PLLLKDET_OUT                      : out  std_logic;
    TILE2_REFCLKOUT_OUT                     : out  std_logic;
    TILE2_RESETDONE0_OUT                    : out  std_logic;
    TILE2_RESETDONE1_OUT                    : out  std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TILE2_TXDATA0_IN                        : in   std_logic_vector(19 downto 0);
    TILE2_TXDATA1_IN                        : in   std_logic_vector(19 downto 0);
    TILE2_TXUSRCLK0_IN                      : in   std_logic;
    TILE2_TXUSRCLK1_IN                      : in   std_logic;
    TILE2_TXUSRCLK20_IN                     : in   std_logic;
    TILE2_TXUSRCLK21_IN                     : in   std_logic;
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    TILE2_TXN0_OUT                          : out  std_logic;
    TILE2_TXN1_OUT                          : out  std_logic;
    TILE2_TXP0_OUT                          : out  std_logic;
    TILE2_TXP1_OUT                          : out  std_logic


);
end component;


component MGT_USRCLK_SOURCE 
generic
(
    FREQUENCY_MODE   : string   := "LOW";    
    PERFORMANCE_MODE : string   := "MAX_SPEED"    
);
port
(
    DIV1_OUT                : out std_logic;
    DIV2_OUT                : out std_logic;
    DCM_LOCKED_OUT          : out std_logic;
    CLK_IN                  : in  std_logic;
    DCM_RESET_IN            : in  std_logic

);
end component;

component FRAME_GEN 
generic
(
    WORDS_IN_BRAM : integer    :=   256;
    MEM_00       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_01       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_02       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_03       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_04       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_05       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_06       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_07       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_08       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_09       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_10       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_11       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_12       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_13       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_14       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_15       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_16       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_17       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_18       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_19       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_20       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_21       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_22       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_23       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_24       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_25       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_26       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_27       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_28       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_29       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_30       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_31       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_32       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_33       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_34       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_35       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_36       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_37       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_38       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_39       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_00      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_01      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_02      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_03      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_04      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_05      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_06      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_07      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000"
);    
port
(
    -- User Interface
    TX_DATA             : out   std_logic_vector(39 downto 0);
    TX_CHARISK          : out   std_logic_vector(3 downto 0); 

    -- System Interface
    USER_CLK            : in    std_logic;
    SYSTEM_RESET        : in    std_logic
); 
end component;

component FRAME_CHECK 
generic
(
    RX_DATA_WIDTH            : integer := 16;
    USE_COMMA                : integer := 1;
    NONE_MSB_FIRST_DEC       : integer := 0;
    COMMA_DOUBLE_DEC         : integer := 0;
    CHANBOND_SEQ_LEN         : integer := 1;
    WORDS_IN_BRAM            : integer := 256;
    CONFIG_INDEPENDENT_LANES : integer := 0;
    START_OF_PACKET_CHAR     : std_logic_vector := x"55fb";
    COMMA_DOUBLE_CHAR        : std_logic_vector := x"f628";
    MEM_00       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_01       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_02       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_03       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_04       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_05       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_06       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_07       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_08       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_09       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_10       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_11       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_12       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_13       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_14       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_15       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_16       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_17       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_18       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_19       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_20       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_21       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_22       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_23       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_24       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_25       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_26       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_27       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_28       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_29       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_30       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_31       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_32       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_33       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_34       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_35       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_36       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_37       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_38       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_39       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_00      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_01      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_02      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_03      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_04      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_05      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_06      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_07      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000"
);
port
(
    -- User Interface
    RX_DATA                  : in  std_logic_vector((RX_DATA_WIDTH-1) downto 0); 
    RX_ENMCOMMA_ALIGN        : out std_logic;
    RX_ENPCOMMA_ALIGN        : out std_logic;
    RX_ENCHAN_SYNC           : out std_logic; 
    RX_CHANBOND_SEQ          : in  std_logic; 

    -- Control Interface
    INC_IN                   : in std_logic; 
    INC_OUT                  : out std_logic; 
    PATTERN_MATCH_N          : out std_logic;
    RESET_ON_ERROR           : in std_logic; 
    
    -- Error Monitoring
    ERROR_COUNT              : out std_logic_vector(7 downto 0);

    -- System Interface
    USER_CLK                 : in std_logic;
    SYSTEM_RESET             : in std_logic
  
);
end component;

component MGT_USRCLK_SOURCE_PLL 
generic
(
    MULT                 : integer          := 2;
    DIVIDE               : integer          := 2;    
    CLK_PERIOD           : real             := 10.0;    
    OUT0_DIVIDE          : integer          := 2;
    OUT1_DIVIDE          : integer          := 2;
    OUT2_DIVIDE          : integer          := 2;
    OUT3_DIVIDE          : integer          := 2;
    SIMULATION_P         : integer          := 1;
    LOCK_WAIT_COUNT      : std_logic_vector := "1000001000110101"  
);
port
( 
    CLK0_OUT                : out std_logic;
    CLK1_OUT                : out std_logic;
    CLK2_OUT                : out std_logic;
    CLK3_OUT                : out std_logic;
    CLK_IN                  : in  std_logic;
    PLL_LOCKED_OUT          : out std_logic;
    PLL_RESET_IN            : in  std_logic
);
end component;






-- Chipscope modules
attribute syn_black_box                : boolean;
attribute syn_noprune                  : boolean;


component shared_vio
port
(
    control                 : in  std_logic_vector(35 downto 0);
    async_in                : in  std_logic_vector(31 downto 0);
    async_out               : out std_logic_vector(31 downto 0)
);
end component;
attribute syn_black_box of shared_vio : component is TRUE;
attribute syn_noprune of shared_vio   : component is TRUE;

component icon
port
(
    control0                : out std_logic_vector(35 downto 0);
    control1                : out std_logic_vector(35 downto 0);
    control2                : out std_logic_vector(35 downto 0);
    control3                : out std_logic_vector(35 downto 0);
    control4                : out std_logic_vector(35 downto 0);
    control5                : out std_logic_vector(35 downto 0);
    control6                : out std_logic_vector(35 downto 0));
end component;


attribute syn_black_box of icon : component is TRUE;
attribute syn_noprune of icon   : component is TRUE;


component ila
port
(
    control                 : in  std_logic_vector(35 downto 0);
    clk                     : in  std_logic;
    trig0                   : in  std_logic_vector(84 downto 0)
);
end component;
attribute syn_black_box of ila : component is TRUE;
attribute syn_noprune of ila   : component is TRUE;


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

    
--************************** Register Declarations ****************************

    signal   tile0_tx_resetdone0_r           : std_logic;
    signal   tile0_tx_resetdone0_r2          : std_logic;
    signal   tile0_rx_resetdone0_r           : std_logic;
    signal   tile0_rx_resetdone0_r2          : std_logic;
    signal   tile0_tx_resetdone1_r           : std_logic;
    signal   tile0_tx_resetdone1_r2          : std_logic;
    signal   tile0_rx_resetdone1_r           : std_logic;
    signal   tile0_rx_resetdone1_r2          : std_logic;
    signal   tile1_tx_resetdone0_r           : std_logic;
    signal   tile1_tx_resetdone0_r2          : std_logic;
    signal   tile1_rx_resetdone0_r           : std_logic;
    signal   tile1_rx_resetdone0_r2          : std_logic;
    signal   tile1_tx_resetdone1_r           : std_logic;
    signal   tile1_tx_resetdone1_r2          : std_logic;
    signal   tile1_rx_resetdone1_r           : std_logic;
    signal   tile1_rx_resetdone1_r2          : std_logic;
    signal   tile2_tx_resetdone0_r           : std_logic;
    signal   tile2_tx_resetdone0_r2          : std_logic;
    signal   tile2_rx_resetdone0_r           : std_logic;
    signal   tile2_rx_resetdone0_r2          : std_logic;
    signal   tile2_tx_resetdone1_r           : std_logic;
    signal   tile2_tx_resetdone1_r2          : std_logic;
    signal   tile2_rx_resetdone1_r           : std_logic;
    signal   tile2_rx_resetdone1_r2          : std_logic;
    signal   async_mux0_sel_i                : std_logic_vector(1 downto 0);
    signal   not_async_mux0_sel_i            : std_logic_vector(1 downto 0);
    signal   async_mux1_sel_i                : std_logic_vector(1 downto 0);
    signal   not_async_mux1_sel_i            : std_logic_vector(1 downto 0);
  

--**************************** Wire Declarations ******************************

    -------------------------- MGT Wrapper Wires ------------------------------
    
    --________________________________________________________________________
    --________________________________________________________________________
    --TILE0   (X0Y3)

    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    signal  tile0_rxchariscomma0_i          : std_logic_vector(1 downto 0);
    signal  tile0_rxchariscomma1_i          : std_logic_vector(1 downto 0);
    signal  tile0_rxdisperr0_i              : std_logic_vector(1 downto 0);
    signal  tile0_rxdisperr1_i              : std_logic_vector(1 downto 0);
    signal  tile0_rxnotintable0_i           : std_logic_vector(1 downto 0);
    signal  tile0_rxnotintable1_i           : std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  tile0_rxbyteisaligned0_i        : std_logic;
    signal  tile0_rxbyteisaligned1_i        : std_logic;
    signal  tile0_rxenmcommaalign0_i        : std_logic;
    signal  tile0_rxenmcommaalign1_i        : std_logic;
    signal  tile0_rxenpcommaalign0_i        : std_logic;
    signal  tile0_rxenpcommaalign1_i        : std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    signal  tile0_rxdata0_i                 : std_logic_vector(15 downto 0);
    signal  tile0_rxdata1_i                 : std_logic_vector(15 downto 0);
    signal  tile0_rxrecclk0_i               : std_logic;
    signal  tile0_rxrecclk1_i               : std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    signal  tile0_rxeqmix0_i                : std_logic_vector(1 downto 0);
    signal  tile0_rxeqmix1_i                : std_logic_vector(1 downto 0);
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    signal  tile0_rxpolarity0_i             : std_logic;
    signal  tile0_rxpolarity1_i             : std_logic;
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    signal  tile0_gtxreset_i                : std_logic;
    signal  tile0_plllkdet_i                : std_logic;
    signal  tile0_refclkout_i               : std_logic;
    signal  tile0_resetdone0_i              : std_logic;
    signal  tile0_resetdone1_i              : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  tile0_txdata0_i                 : std_logic_vector(19 downto 0);
    signal  tile0_txdata1_i                 : std_logic_vector(19 downto 0);


    --________________________________________________________________________
    --________________________________________________________________________
    --TILE1   (X0Y4)

    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    signal  tile1_rxchariscomma0_i          : std_logic_vector(1 downto 0);
    signal  tile1_rxchariscomma1_i          : std_logic_vector(1 downto 0);
    signal  tile1_rxdisperr0_i              : std_logic_vector(1 downto 0);
    signal  tile1_rxdisperr1_i              : std_logic_vector(1 downto 0);
    signal  tile1_rxnotintable0_i           : std_logic_vector(1 downto 0);
    signal  tile1_rxnotintable1_i           : std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  tile1_rxbyteisaligned0_i        : std_logic;
    signal  tile1_rxbyteisaligned1_i        : std_logic;
    signal  tile1_rxenmcommaalign0_i        : std_logic;
    signal  tile1_rxenmcommaalign1_i        : std_logic;
    signal  tile1_rxenpcommaalign0_i        : std_logic;
    signal  tile1_rxenpcommaalign1_i        : std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    signal  tile1_rxdata0_i                 : std_logic_vector(15 downto 0);
    signal  tile1_rxdata1_i                 : std_logic_vector(15 downto 0);
    signal  tile1_rxrecclk0_i               : std_logic;
    signal  tile1_rxrecclk1_i               : std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    signal  tile1_rxeqmix0_i                : std_logic_vector(1 downto 0);
    signal  tile1_rxeqmix1_i                : std_logic_vector(1 downto 0);
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    signal  tile1_rxpolarity0_i             : std_logic;
    signal  tile1_rxpolarity1_i             : std_logic;
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    signal  tile1_gtxreset_i                : std_logic;
    signal  tile1_plllkdet_i                : std_logic;
    signal  tile1_refclkout_i               : std_logic;
    signal  tile1_resetdone0_i              : std_logic;
    signal  tile1_resetdone1_i              : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  tile1_txdata0_i                 : std_logic_vector(19 downto 0);
    signal  tile1_txdata1_i                 : std_logic_vector(19 downto 0);


    --________________________________________________________________________
    --________________________________________________________________________
    --TILE2   (X0Y5)

    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    signal  tile2_rxchariscomma0_i          : std_logic_vector(1 downto 0);
    signal  tile2_rxchariscomma1_i          : std_logic_vector(1 downto 0);
    signal  tile2_rxdisperr0_i              : std_logic_vector(1 downto 0);
    signal  tile2_rxdisperr1_i              : std_logic_vector(1 downto 0);
    signal  tile2_rxnotintable0_i           : std_logic_vector(1 downto 0);
    signal  tile2_rxnotintable1_i           : std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  tile2_rxbyteisaligned0_i        : std_logic;
    signal  tile2_rxbyteisaligned1_i        : std_logic;
    signal  tile2_rxenmcommaalign0_i        : std_logic;
    signal  tile2_rxenmcommaalign1_i        : std_logic;
    signal  tile2_rxenpcommaalign0_i        : std_logic;
    signal  tile2_rxenpcommaalign1_i        : std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    signal  tile2_rxdata0_i                 : std_logic_vector(15 downto 0);
    signal  tile2_rxdata1_i                 : std_logic_vector(15 downto 0);
    signal  tile2_rxrecclk0_i               : std_logic;
    signal  tile2_rxrecclk1_i               : std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    signal  tile2_rxeqmix0_i                : std_logic_vector(1 downto 0);
    signal  tile2_rxeqmix1_i                : std_logic_vector(1 downto 0);
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    signal  tile2_rxpolarity0_i             : std_logic;
    signal  tile2_rxpolarity1_i             : std_logic;
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    signal  tile2_gtxreset_i                : std_logic;
    signal  tile2_plllkdet_i                : std_logic;
    signal  tile2_refclkout_i               : std_logic;
    signal  tile2_resetdone0_i              : std_logic;
    signal  tile2_resetdone1_i              : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  tile2_txdata0_i                 : std_logic_vector(19 downto 0);
    signal  tile2_txdata1_i                 : std_logic_vector(19 downto 0);


    ------------------------------- Global Signals -----------------------------
    signal  tile0_tx_system_reset0_c        : std_logic;
    signal  tile0_rx_system_reset0_c        : std_logic;
    signal  tile0_tx_system_reset1_c        : std_logic;
    signal  tile0_rx_system_reset1_c        : std_logic;
    signal  tile1_tx_system_reset0_c        : std_logic;
    signal  tile1_rx_system_reset0_c        : std_logic;
    signal  tile1_tx_system_reset1_c        : std_logic;
    signal  tile1_rx_system_reset1_c        : std_logic;
    signal  tile2_tx_system_reset0_c        : std_logic;
    signal  tile2_rx_system_reset0_c        : std_logic;
    signal  tile2_tx_system_reset1_c        : std_logic;
    signal  tile2_rx_system_reset1_c        : std_logic;
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_ground_vec_i            : std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   : std_logic;
    signal  tied_to_vcc_vec_i               : std_logic_vector(7 downto 0);
    signal  drp_clk_in_i                    : std_logic;
    
    signal  tile0_refclkout_bufg_i          : std_logic;
    
    
    ----------------------------- User Clocks ---------------------------------
    signal  tile0_txusrclk0_i               : std_logic;
    signal  tile0_rxusrclk0_i               : std_logic;
    signal  tile0_rxusrclk1_i               : std_logic;
    signal  tile1_rxusrclk0_i               : std_logic;
    signal  tile1_rxusrclk1_i               : std_logic;
    signal  tile2_rxusrclk0_i               : std_logic;
    signal  tile2_rxusrclk1_i               : std_logic;


    ----------------------- Frame check/gen Module Signals --------------------
    signal  tile0_matchn0_i                 : std_logic;
     
    signal  tile0_txcharisk0_float_i        : std_logic_vector(1 downto 0);
    signal  tile0_txdata0_float_i           : std_logic_vector(19 downto 0);
    
    
    signal  tile0_block_sync0_i             : std_logic;
    signal  tile0_error_count0_i            : std_logic_vector(7 downto 0);
    signal  tile0_frame_check0_reset_i      : std_logic;
    signal  tile0_inc_in0_i                 : std_logic;
    signal  tile0_inc_out0_i                : std_logic;
    signal  tile0_unscrambled_data0_i       : std_logic_vector(15 downto 0);
    signal  tile0_matchn1_i                 : std_logic;
     
    signal  tile0_txcharisk1_float_i        : std_logic_vector(1 downto 0);
    signal  tile0_txdata1_float_i           : std_logic_vector(19 downto 0);
    
    
    signal  tile0_block_sync1_i             : std_logic;
    signal  tile0_error_count1_i            : std_logic_vector(7 downto 0);
    signal  tile0_frame_check1_reset_i      : std_logic;
    signal  tile0_inc_in1_i                 : std_logic;
    signal  tile0_inc_out1_i                : std_logic;
    signal  tile0_unscrambled_data1_i       : std_logic_vector(15 downto 0);

    signal  tile1_matchn0_i                 : std_logic;
     
    signal  tile1_txcharisk0_float_i        : std_logic_vector(1 downto 0);
    signal  tile1_txdata0_float_i           : std_logic_vector(19 downto 0);
    
    
    signal  tile1_block_sync0_i             : std_logic;
    signal  tile1_error_count0_i            : std_logic_vector(7 downto 0);
    signal  tile1_frame_check0_reset_i      : std_logic;
    signal  tile1_inc_in0_i                 : std_logic;
    signal  tile1_inc_out0_i                : std_logic;
    signal  tile1_unscrambled_data0_i       : std_logic_vector(15 downto 0);
    signal  tile1_matchn1_i                 : std_logic;
     
    signal  tile1_txcharisk1_float_i        : std_logic_vector(1 downto 0);
    signal  tile1_txdata1_float_i           : std_logic_vector(19 downto 0);
    
    
    signal  tile1_block_sync1_i             : std_logic;
    signal  tile1_error_count1_i            : std_logic_vector(7 downto 0);
    signal  tile1_frame_check1_reset_i      : std_logic;
    signal  tile1_inc_in1_i                 : std_logic;
    signal  tile1_inc_out1_i                : std_logic;
    signal  tile1_unscrambled_data1_i       : std_logic_vector(15 downto 0);

    signal  tile2_refclk_i                  : std_logic;
    signal  tile2_matchn0_i                 : std_logic;
     
    signal  tile2_txcharisk0_float_i        : std_logic_vector(1 downto 0);
    signal  tile2_txdata0_float_i           : std_logic_vector(19 downto 0);
    
    
    signal  tile2_block_sync0_i             : std_logic;
    signal  tile2_error_count0_i            : std_logic_vector(7 downto 0);
    signal  tile2_frame_check0_reset_i      : std_logic;
    signal  tile2_inc_in0_i                 : std_logic;
    signal  tile2_inc_out0_i                : std_logic;
    signal  tile2_unscrambled_data0_i       : std_logic_vector(15 downto 0);
    signal  tile2_matchn1_i                 : std_logic;
     
    signal  tile2_txcharisk1_float_i        : std_logic_vector(1 downto 0);
    signal  tile2_txdata1_float_i           : std_logic_vector(19 downto 0);
    
    
    signal  tile2_block_sync1_i             : std_logic;
    signal  tile2_error_count1_i            : std_logic_vector(7 downto 0);
    signal  tile2_frame_check1_reset_i      : std_logic;
    signal  tile2_inc_in1_i                 : std_logic;
    signal  tile2_inc_out1_i                : std_logic;
    signal  tile2_unscrambled_data1_i       : std_logic_vector(15 downto 0);

    signal  reset_on_data_error_i           : std_logic;


    ----------------------- Chipscope Signals ---------------------------------

    signal  shared_vio_control_i            : std_logic_vector(35 downto 0);
    signal  tx_data_vio_control0_i          : std_logic_vector(35 downto 0);
    signal  tx_data_vio_control1_i          : std_logic_vector(35 downto 0);
    signal  rx_data_vio_control0_i          : std_logic_vector(35 downto 0);
    signal  rx_data_vio_control1_i          : std_logic_vector(35 downto 0);
    signal  ila_control0_i                  : std_logic_vector(35 downto 0);
    signal  ila_control1_i                  : std_logic_vector(35 downto 0);
    signal  shared_vio_in_i                 : std_logic_vector(31 downto 0);
    signal  shared_vio_out_i                : std_logic_vector(31 downto 0);
    signal  tx_data_vio_in0_i               : std_logic_vector(31 downto 0);
    signal  tx_data_vio_out0_i              : std_logic_vector(31 downto 0);
    signal  tx_data_vio_in1_i               : std_logic_vector(31 downto 0);
    signal  tx_data_vio_out1_i              : std_logic_vector(31 downto 0);
    signal  rx_data_vio_in0_i               : std_logic_vector(31 downto 0);
    signal  rx_data_vio_out0_i              : std_logic_vector(31 downto 0);
    signal  rx_data_vio_in1_i               : std_logic_vector(31 downto 0);
    signal  rx_data_vio_out1_i              : std_logic_vector(31 downto 0);
    signal  ila_in0_i                       : std_logic_vector(84 downto 0);
    signal  ila_in1_i                       : std_logic_vector(84 downto 0);

    signal  tile0_tx_data_vio_in0_i         : std_logic_vector(31 downto 0);
    signal  tile0_tx_data_vio_out0_i        : std_logic_vector(31 downto 0);
    signal  tile0_tx_data_vio_in1_i         : std_logic_vector(31 downto 0);
    signal  tile0_tx_data_vio_out1_i        : std_logic_vector(31 downto 0);
    signal  tile0_rx_data_vio_in0_i         : std_logic_vector(31 downto 0);
    signal  tile0_rx_data_vio_out0_i        : std_logic_vector(31 downto 0);
    signal  tile0_rx_data_vio_in1_i         : std_logic_vector(31 downto 0);
    signal  tile0_rx_data_vio_out1_i        : std_logic_vector(31 downto 0);
    signal  tile0_ila_in0_i                 : std_logic_vector(84 downto 0);
    signal  tile0_ila_in1_i                 : std_logic_vector(84 downto 0);

    signal  tile1_tx_data_vio_in0_i         : std_logic_vector(31 downto 0);
    signal  tile1_tx_data_vio_out0_i        : std_logic_vector(31 downto 0);
    signal  tile1_tx_data_vio_in1_i         : std_logic_vector(31 downto 0);
    signal  tile1_tx_data_vio_out1_i        : std_logic_vector(31 downto 0);
    signal  tile1_rx_data_vio_in0_i         : std_logic_vector(31 downto 0);
    signal  tile1_rx_data_vio_out0_i        : std_logic_vector(31 downto 0);
    signal  tile1_rx_data_vio_in1_i         : std_logic_vector(31 downto 0);
    signal  tile1_rx_data_vio_out1_i        : std_logic_vector(31 downto 0);
    signal  tile1_ila_in0_i                 : std_logic_vector(84 downto 0);
    signal  tile1_ila_in1_i                 : std_logic_vector(84 downto 0);

    signal  tile2_tx_data_vio_in0_i         : std_logic_vector(31 downto 0);
    signal  tile2_tx_data_vio_out0_i        : std_logic_vector(31 downto 0);
    signal  tile2_tx_data_vio_in1_i         : std_logic_vector(31 downto 0);
    signal  tile2_tx_data_vio_out1_i        : std_logic_vector(31 downto 0);
    signal  tile2_rx_data_vio_in0_i         : std_logic_vector(31 downto 0);
    signal  tile2_rx_data_vio_out0_i        : std_logic_vector(31 downto 0);
    signal  tile2_rx_data_vio_in1_i         : std_logic_vector(31 downto 0);
    signal  tile2_rx_data_vio_out1_i        : std_logic_vector(31 downto 0);
    signal  tile2_ila_in0_i                 : std_logic_vector(84 downto 0);
    signal  tile2_ila_in1_i                 : std_logic_vector(84 downto 0);


    signal  gtxreset_i                      : std_logic;
    signal  mux_sel_i                       : std_logic_vector(1 downto 0);
    signal  not_mux_sel_i                   : std_logic_vector(1 downto 0);    
    signal  user_tx_reset_i                 : std_logic;
    signal  user_rx_reset_i                 : std_logic;
    signal  ila_clk0_i                      : std_logic;
    signal  ila_clk1_i                      : std_logic;
    signal ila_clk0_mux_out0_i             : std_logic;
    signal ila_clk1_mux_out0_i             : std_logic;


--**************************** Main Body of Code *******************************
begin

    --  Static signal Assigments
    tied_to_ground_i                        <= '0';
    tied_to_ground_vec_i                    <= x"0000000000000000";
    tied_to_vcc_i                           <= '1';
    tied_to_vcc_vec_i                       <= x"ff";


    




    -----------------------Dedicated GTX Reference Clock Inputs ---------------
    -- The dedicated reference clock inputs you selected in the GUI are implemented using
    -- IBUFDS instances.
    --
    -- In the UCF file for this example design, you will see that each of
    -- these IBUFDS instances has been LOCed to a particular set of pins. By LOCing to these
    -- locations, we tell the tools to use the dedicated input buffers to the GTX reference
    -- clock network, rather than general purpose IOs. To select other pins, consult the 
    -- Implementation chapter of UG196, or rerun the wizard.
    --
    -- This network is the highest performace (lowest jitter) option for providing clocks
    -- to the GTX transceivers.
    
    tile2_refclk_ibufds_i : IBUFDS
    port map
    (
        O                               =>      tile2_refclk_i,
        I                               =>      TILE2_REFCLK_PAD_P_IN,
        IB                              =>      TILE2_REFCLK_PAD_N_IN
    );






    ----------------------------------- User Clocks ---------------------------
    
    -- The clock resources in this section were added based on userclk source selections on
    -- the Latency, Buffering, and Clocking page of the GUI. A few notes about user clocks:
    -- * The userclk and userclk2 for each GTX datapath (TX and RX) must be phase aligned to 
    --   avoid data errors in the fabric interface whenever the datapath is wider than 10 bits
    -- * To minimize clock resources, you can share clocks between GTXs. GTXs using the same frequency
    --   or multiples of the same frequency can be accomadated using DCMs and PLLs. Use caution when
    --   using RXRECCLK as a clock source, however - these clocks can typically only be shared if all
    --   the channels using the clock are receiving data from TX channels that share a reference clock 
    --   source with each other.

    refclkout_bufg0_i : BUFG
    port map
    (
        I                               =>      tile0_refclkout_i,
        O                               =>      tile0_txusrclk0_i
    );


    rxrecclk_bufg1_i : BUFG
    port map
    (
        I                               =>      tile0_rxrecclk0_i,
        O                               =>      tile0_rxusrclk0_i
    );


    rxrecclk_bufg2_i : BUFG
    port map
    (
        I                               =>      tile0_rxrecclk1_i,
        O                               =>      tile0_rxusrclk1_i
    );


    rxrecclk_bufg3_i : BUFG
    port map
    (
        I                               =>      tile1_rxrecclk0_i,
        O                               =>      tile1_rxusrclk0_i
    );


    rxrecclk_bufg4_i : BUFG
    port map
    (
        I                               =>      tile1_rxrecclk1_i,
        O                               =>      tile1_rxusrclk1_i
    );


    rxrecclk_bufg5_i : BUFG
    port map
    (
        I                               =>      tile2_rxrecclk0_i,
        O                               =>      tile2_rxusrclk0_i
    );


    rxrecclk_bufg6_i : BUFG
    port map
    (
        I                               =>      tile2_rxrecclk1_i,
        O                               =>      tile2_rxusrclk1_i
    );






    ----------------------------- The GTX Wrapper -----------------------------
    
    -- Use the instantiation template in the examples directory to add the GTX wrapper to your design.
    -- In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    -- checker. The GTXs will reset, then attempt to align and transmit data. If channel bonding is 
    -- enabled, bonding should occur after alignment.


    -- Wire all PLLLKDET signals to the top level as output ports
    TILE0_PLLLKDET_OUT                      <= tile0_plllkdet_i;
    TILE1_PLLLKDET_OUT                      <= tile1_plllkdet_i;
    TILE2_PLLLKDET_OUT                      <= tile2_plllkdet_i;



    gtx_i : GTX
    generic map
    (
        WRAPPER_SIM_MODE                =>      EXAMPLE_SIM_MODE,
        WRAPPER_SIM_GTXRESET_SPEEDUP    =>      EXAMPLE_SIM_GTXRESET_SPEEDUP,
        WRAPPER_SIM_PLL_PERDIV2         =>      EXAMPLE_SIM_PLL_PERDIV2
    )
    port map
    (
    
 
 
 
 
 
 
 
 
        --_____________________________________________________________________
        --_____________________________________________________________________
        --TILE0  (X0Y3)

        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        TILE0_RXCHARISCOMMA0_OUT        =>      tile0_rxchariscomma0_i,
        TILE0_RXCHARISCOMMA1_OUT        =>      tile0_rxchariscomma1_i,
        TILE0_RXDISPERR0_OUT            =>      tile0_rxdisperr0_i,
        TILE0_RXDISPERR1_OUT            =>      tile0_rxdisperr1_i,
        TILE0_RXNOTINTABLE0_OUT         =>      tile0_rxnotintable0_i,
        TILE0_RXNOTINTABLE1_OUT         =>      tile0_rxnotintable1_i,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        TILE0_RXBYTEISALIGNED0_OUT      =>      tile0_rxbyteisaligned0_i,
        TILE0_RXBYTEISALIGNED1_OUT      =>      tile0_rxbyteisaligned1_i,
        TILE0_RXENMCOMMAALIGN0_IN       =>      tile0_rxenmcommaalign0_i,
        TILE0_RXENMCOMMAALIGN1_IN       =>      tile0_rxenmcommaalign1_i,
        TILE0_RXENPCOMMAALIGN0_IN       =>      tile0_rxenpcommaalign0_i,
        TILE0_RXENPCOMMAALIGN1_IN       =>      tile0_rxenpcommaalign1_i,
        ------------------- Receive Ports - RX Data Path interface -----------------
        TILE0_RXDATA0_OUT               =>      tile0_rxdata0_i,
        TILE0_RXDATA1_OUT               =>      tile0_rxdata1_i,
        TILE0_RXRECCLK0_OUT             =>      tile0_rxrecclk0_i,
        TILE0_RXRECCLK1_OUT             =>      tile0_rxrecclk1_i,
        TILE0_RXUSRCLK0_IN              =>      tile0_rxusrclk0_i,
        TILE0_RXUSRCLK1_IN              =>      tile0_rxusrclk1_i,
        TILE0_RXUSRCLK20_IN             =>      tile0_rxusrclk0_i,
        TILE0_RXUSRCLK21_IN             =>      tile0_rxusrclk1_i,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        TILE0_RXEQMIX0_IN               =>      tile0_rxeqmix0_i,
        TILE0_RXEQMIX1_IN               =>      tile0_rxeqmix1_i,
        TILE0_RXN0_IN                   =>      RXN_IN(0),
        TILE0_RXN1_IN                   =>      RXN_IN(1),
        TILE0_RXP0_IN                   =>      RXP_IN(0),
        TILE0_RXP1_IN                   =>      RXP_IN(1),
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        TILE0_RXPOLARITY0_IN            =>      tile0_rxpolarity0_i,
        TILE0_RXPOLARITY1_IN            =>      tile0_rxpolarity1_i,
        --------------------- Shared Ports - Tile and PLL Ports --------------------
        TILE0_CLKIN_IN                  =>      tile2_refclk_i,
        TILE0_GTXRESET_IN               =>      tile0_gtxreset_i,
        TILE0_PLLLKDET_OUT              =>      tile0_plllkdet_i,
        TILE0_REFCLKOUT_OUT             =>      tile0_refclkout_i,
        TILE0_RESETDONE0_OUT            =>      tile0_resetdone0_i,
        TILE0_RESETDONE1_OUT            =>      tile0_resetdone1_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TILE0_TXDATA0_IN                =>      tile0_txdata0_i,
        TILE0_TXDATA1_IN                =>      tile0_txdata1_i,
        TILE0_TXUSRCLK0_IN              =>      tile0_txusrclk0_i,
        TILE0_TXUSRCLK1_IN              =>      tile0_txusrclk0_i,
        TILE0_TXUSRCLK20_IN             =>      tile0_txusrclk0_i,
        TILE0_TXUSRCLK21_IN             =>      tile0_txusrclk0_i,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TILE0_TXN0_OUT                  =>      TXN_OUT(0),
        TILE0_TXN1_OUT                  =>      TXN_OUT(1),
        TILE0_TXP0_OUT                  =>      TXP_OUT(0),
        TILE0_TXP1_OUT                  =>      TXP_OUT(1),


    
 
 
 
 
 
 
 
 
        --_____________________________________________________________________
        --_____________________________________________________________________
        --TILE1  (X0Y4)

        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        TILE1_RXCHARISCOMMA0_OUT        =>      tile1_rxchariscomma0_i,
        TILE1_RXCHARISCOMMA1_OUT        =>      tile1_rxchariscomma1_i,
        TILE1_RXDISPERR0_OUT            =>      tile1_rxdisperr0_i,
        TILE1_RXDISPERR1_OUT            =>      tile1_rxdisperr1_i,
        TILE1_RXNOTINTABLE0_OUT         =>      tile1_rxnotintable0_i,
        TILE1_RXNOTINTABLE1_OUT         =>      tile1_rxnotintable1_i,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        TILE1_RXBYTEISALIGNED0_OUT      =>      tile1_rxbyteisaligned0_i,
        TILE1_RXBYTEISALIGNED1_OUT      =>      tile1_rxbyteisaligned1_i,
        TILE1_RXENMCOMMAALIGN0_IN       =>      tile1_rxenmcommaalign0_i,
        TILE1_RXENMCOMMAALIGN1_IN       =>      tile1_rxenmcommaalign1_i,
        TILE1_RXENPCOMMAALIGN0_IN       =>      tile1_rxenpcommaalign0_i,
        TILE1_RXENPCOMMAALIGN1_IN       =>      tile1_rxenpcommaalign1_i,
        ------------------- Receive Ports - RX Data Path interface -----------------
        TILE1_RXDATA0_OUT               =>      tile1_rxdata0_i,
        TILE1_RXDATA1_OUT               =>      tile1_rxdata1_i,
        TILE1_RXRECCLK0_OUT             =>      tile1_rxrecclk0_i,
        TILE1_RXRECCLK1_OUT             =>      tile1_rxrecclk1_i,
        TILE1_RXUSRCLK0_IN              =>      tile1_rxusrclk0_i,
        TILE1_RXUSRCLK1_IN              =>      tile1_rxusrclk1_i,
        TILE1_RXUSRCLK20_IN             =>      tile1_rxusrclk0_i,
        TILE1_RXUSRCLK21_IN             =>      tile1_rxusrclk1_i,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        TILE1_RXEQMIX0_IN               =>      tile1_rxeqmix0_i,
        TILE1_RXEQMIX1_IN               =>      tile1_rxeqmix1_i,
        TILE1_RXN0_IN                   =>      RXN_IN(2),
        TILE1_RXN1_IN                   =>      RXN_IN(3),
        TILE1_RXP0_IN                   =>      RXP_IN(2),
        TILE1_RXP1_IN                   =>      RXP_IN(3),
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        TILE1_RXPOLARITY0_IN            =>      tile1_rxpolarity0_i,
        TILE1_RXPOLARITY1_IN            =>      tile1_rxpolarity1_i,
        --------------------- Shared Ports - Tile and PLL Ports --------------------
        TILE1_CLKIN_IN                  =>      tile2_refclk_i,
        TILE1_GTXRESET_IN               =>      tile1_gtxreset_i,
        TILE1_PLLLKDET_OUT              =>      tile1_plllkdet_i,
        TILE1_REFCLKOUT_OUT             =>      tile1_refclkout_i,
        TILE1_RESETDONE0_OUT            =>      tile1_resetdone0_i,
        TILE1_RESETDONE1_OUT            =>      tile1_resetdone1_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TILE1_TXDATA0_IN                =>      tile1_txdata0_i,
        TILE1_TXDATA1_IN                =>      tile1_txdata1_i,
        TILE1_TXUSRCLK0_IN              =>      tile0_txusrclk0_i,
        TILE1_TXUSRCLK1_IN              =>      tile0_txusrclk0_i,
        TILE1_TXUSRCLK20_IN             =>      tile0_txusrclk0_i,
        TILE1_TXUSRCLK21_IN             =>      tile0_txusrclk0_i,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TILE1_TXN0_OUT                  =>      TXN_OUT(2),
        TILE1_TXN1_OUT                  =>      TXN_OUT(3),
        TILE1_TXP0_OUT                  =>      TXP_OUT(2),
        TILE1_TXP1_OUT                  =>      TXP_OUT(3),


    
 
 
 
 
 
 
 
 
        --_____________________________________________________________________
        --_____________________________________________________________________
        --TILE2  (X0Y5)

        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        TILE2_RXCHARISCOMMA0_OUT        =>      tile2_rxchariscomma0_i,
        TILE2_RXCHARISCOMMA1_OUT        =>      tile2_rxchariscomma1_i,
        TILE2_RXDISPERR0_OUT            =>      tile2_rxdisperr0_i,
        TILE2_RXDISPERR1_OUT            =>      tile2_rxdisperr1_i,
        TILE2_RXNOTINTABLE0_OUT         =>      tile2_rxnotintable0_i,
        TILE2_RXNOTINTABLE1_OUT         =>      tile2_rxnotintable1_i,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        TILE2_RXBYTEISALIGNED0_OUT      =>      tile2_rxbyteisaligned0_i,
        TILE2_RXBYTEISALIGNED1_OUT      =>      tile2_rxbyteisaligned1_i,
        TILE2_RXENMCOMMAALIGN0_IN       =>      tile2_rxenmcommaalign0_i,
        TILE2_RXENMCOMMAALIGN1_IN       =>      tile2_rxenmcommaalign1_i,
        TILE2_RXENPCOMMAALIGN0_IN       =>      tile2_rxenpcommaalign0_i,
        TILE2_RXENPCOMMAALIGN1_IN       =>      tile2_rxenpcommaalign1_i,
        ------------------- Receive Ports - RX Data Path interface -----------------
        TILE2_RXDATA0_OUT               =>      tile2_rxdata0_i,
        TILE2_RXDATA1_OUT               =>      tile2_rxdata1_i,
        TILE2_RXRECCLK0_OUT             =>      tile2_rxrecclk0_i,
        TILE2_RXRECCLK1_OUT             =>      tile2_rxrecclk1_i,
        TILE2_RXUSRCLK0_IN              =>      tile2_rxusrclk0_i,
        TILE2_RXUSRCLK1_IN              =>      tile2_rxusrclk1_i,
        TILE2_RXUSRCLK20_IN             =>      tile2_rxusrclk0_i,
        TILE2_RXUSRCLK21_IN             =>      tile2_rxusrclk1_i,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        TILE2_RXEQMIX0_IN               =>      tile2_rxeqmix0_i,
        TILE2_RXEQMIX1_IN               =>      tile2_rxeqmix1_i,
        TILE2_RXN0_IN                   =>      RXN_IN(4),
        TILE2_RXN1_IN                   =>      RXN_IN(5),
        TILE2_RXP0_IN                   =>      RXP_IN(4),
        TILE2_RXP1_IN                   =>      RXP_IN(5),
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        TILE2_RXPOLARITY0_IN            =>      tile2_rxpolarity0_i,
        TILE2_RXPOLARITY1_IN            =>      tile2_rxpolarity1_i,
        --------------------- Shared Ports - Tile and PLL Ports --------------------
        TILE2_CLKIN_IN                  =>      tile2_refclk_i,
        TILE2_GTXRESET_IN               =>      tile2_gtxreset_i,
        TILE2_PLLLKDET_OUT              =>      tile2_plllkdet_i,
        TILE2_REFCLKOUT_OUT             =>      tile2_refclkout_i,
        TILE2_RESETDONE0_OUT            =>      tile2_resetdone0_i,
        TILE2_RESETDONE1_OUT            =>      tile2_resetdone1_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TILE2_TXDATA0_IN                =>      tile2_txdata0_i,
        TILE2_TXDATA1_IN                =>      tile2_txdata1_i,
        TILE2_TXUSRCLK0_IN              =>      tile0_txusrclk0_i,
        TILE2_TXUSRCLK1_IN              =>      tile0_txusrclk0_i,
        TILE2_TXUSRCLK20_IN             =>      tile0_txusrclk0_i,
        TILE2_TXUSRCLK21_IN             =>      tile0_txusrclk0_i,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TILE2_TXN0_OUT                  =>      TXN_OUT(4),
        TILE2_TXN1_OUT                  =>      TXN_OUT(5),
        TILE2_TXP0_OUT                  =>      TXP_OUT(4),
        TILE2_TXP1_OUT                  =>      TXP_OUT(5)


    );







    -------------------------- User Module Resets -----------------------------
    -- All the User Modules i.e. FRAME_GEN, FRAME_CHECK and the sync modules
    -- are held in reset till the RESETDONE goes high. 
    -- The RESETDONE is registered a couple of times on USRCLK2 and connected 
    -- to the reset of the modules
    
    process( tile0_rxusrclk0_i,tile0_resetdone0_i)
    begin
        if(tile0_resetdone0_i = '0') then
            tile0_rx_resetdone0_r  <= '0'   after DLY;
            tile0_rx_resetdone0_r2 <= '0'   after DLY;
        elsif(tile0_rxusrclk0_i'event and tile0_rxusrclk0_i = '1') then
            tile0_rx_resetdone0_r  <= tile0_resetdone0_i   after DLY;
            tile0_rx_resetdone0_r2 <= tile0_rx_resetdone0_r   after DLY;
        end if;
    end process;
    process( tile0_txusrclk0_i,tile0_resetdone0_i)
    begin
        if(tile0_resetdone0_i = '0') then
            tile0_tx_resetdone0_r  <= '0'   after DLY;
            tile0_tx_resetdone0_r2 <= '0'   after DLY;
        elsif(tile0_txusrclk0_i'event and tile0_txusrclk0_i = '1') then
            tile0_tx_resetdone0_r  <= tile0_resetdone0_i   after DLY;
            tile0_tx_resetdone0_r2 <= tile0_tx_resetdone0_r   after DLY;
        end if;
    end process;
    process( tile0_rxusrclk1_i,tile0_resetdone1_i)
    begin
        if(tile0_resetdone1_i = '0') then
            tile0_rx_resetdone1_r  <= '0'   after DLY;
            tile0_rx_resetdone1_r2 <= '0'   after DLY;
        elsif(tile0_rxusrclk1_i'event and tile0_rxusrclk1_i = '1') then
            tile0_rx_resetdone1_r  <= tile0_resetdone1_i   after DLY;
            tile0_rx_resetdone1_r2 <= tile0_rx_resetdone1_r   after DLY;
        end if;
    end process;
    process( tile0_txusrclk0_i,tile0_resetdone1_i)
    begin
        if(tile0_resetdone1_i = '0') then
            tile0_tx_resetdone1_r  <= '0'   after DLY;
            tile0_tx_resetdone1_r2 <= '0'   after DLY;
        elsif(tile0_txusrclk0_i'event and tile0_txusrclk0_i = '1') then
            tile0_tx_resetdone1_r  <= tile0_resetdone1_i   after DLY;
            tile0_tx_resetdone1_r2 <= tile0_tx_resetdone1_r   after DLY;
        end if;
    end process;
    process( tile1_rxusrclk0_i,tile1_resetdone0_i)
    begin
        if(tile1_resetdone0_i = '0') then
            tile1_rx_resetdone0_r  <= '0'   after DLY;
            tile1_rx_resetdone0_r2 <= '0'   after DLY;
        elsif(tile1_rxusrclk0_i'event and tile1_rxusrclk0_i = '1') then
            tile1_rx_resetdone0_r  <= tile1_resetdone0_i   after DLY;
            tile1_rx_resetdone0_r2 <= tile1_rx_resetdone0_r   after DLY;
        end if;
    end process;
    process( tile0_txusrclk0_i,tile1_resetdone0_i)
    begin
        if(tile1_resetdone0_i = '0') then
            tile1_tx_resetdone0_r  <= '0'   after DLY;
            tile1_tx_resetdone0_r2 <= '0'   after DLY;
        elsif(tile0_txusrclk0_i'event and tile0_txusrclk0_i = '1') then
            tile1_tx_resetdone0_r  <= tile1_resetdone0_i   after DLY;
            tile1_tx_resetdone0_r2 <= tile1_tx_resetdone0_r   after DLY;
        end if;
    end process;
    process( tile1_rxusrclk1_i,tile1_resetdone1_i)
    begin
        if(tile1_resetdone1_i = '0') then
            tile1_rx_resetdone1_r  <= '0'   after DLY;
            tile1_rx_resetdone1_r2 <= '0'   after DLY;
        elsif(tile1_rxusrclk1_i'event and tile1_rxusrclk1_i = '1') then
            tile1_rx_resetdone1_r  <= tile1_resetdone1_i   after DLY;
            tile1_rx_resetdone1_r2 <= tile1_rx_resetdone1_r   after DLY;
        end if;
    end process;
    process( tile0_txusrclk0_i,tile1_resetdone1_i)
    begin
        if(tile1_resetdone1_i = '0') then
            tile1_tx_resetdone1_r  <= '0'   after DLY;
            tile1_tx_resetdone1_r2 <= '0'   after DLY;
        elsif(tile0_txusrclk0_i'event and tile0_txusrclk0_i = '1') then
            tile1_tx_resetdone1_r  <= tile1_resetdone1_i   after DLY;
            tile1_tx_resetdone1_r2 <= tile1_tx_resetdone1_r   after DLY;
        end if;
    end process;
    process( tile2_rxusrclk0_i,tile2_resetdone0_i)
    begin
        if(tile2_resetdone0_i = '0') then
            tile2_rx_resetdone0_r  <= '0'   after DLY;
            tile2_rx_resetdone0_r2 <= '0'   after DLY;
        elsif(tile2_rxusrclk0_i'event and tile2_rxusrclk0_i = '1') then
            tile2_rx_resetdone0_r  <= tile2_resetdone0_i   after DLY;
            tile2_rx_resetdone0_r2 <= tile2_rx_resetdone0_r   after DLY;
        end if;
    end process;
    process( tile0_txusrclk0_i,tile2_resetdone0_i)
    begin
        if(tile2_resetdone0_i = '0') then
            tile2_tx_resetdone0_r  <= '0'   after DLY;
            tile2_tx_resetdone0_r2 <= '0'   after DLY;
        elsif(tile0_txusrclk0_i'event and tile0_txusrclk0_i = '1') then
            tile2_tx_resetdone0_r  <= tile2_resetdone0_i   after DLY;
            tile2_tx_resetdone0_r2 <= tile2_tx_resetdone0_r   after DLY;
        end if;
    end process;
    process( tile2_rxusrclk1_i,tile2_resetdone1_i)
    begin
        if(tile2_resetdone1_i = '0') then
            tile2_rx_resetdone1_r  <= '0'   after DLY;
            tile2_rx_resetdone1_r2 <= '0'   after DLY;
        elsif(tile2_rxusrclk1_i'event and tile2_rxusrclk1_i = '1') then
            tile2_rx_resetdone1_r  <= tile2_resetdone1_i   after DLY;
            tile2_rx_resetdone1_r2 <= tile2_rx_resetdone1_r   after DLY;
        end if;
    end process;
    process( tile0_txusrclk0_i,tile2_resetdone1_i)
    begin
        if(tile2_resetdone1_i = '0') then
            tile2_tx_resetdone1_r  <= '0'   after DLY;
            tile2_tx_resetdone1_r2 <= '0'   after DLY;
        elsif(tile0_txusrclk0_i'event and tile0_txusrclk0_i = '1') then
            tile2_tx_resetdone1_r  <= tile2_resetdone1_i   after DLY;
            tile2_tx_resetdone1_r2 <= tile2_tx_resetdone1_r   after DLY;
        end if;
    end process;

    



    ------------------------------ Frame Generators ---------------------------
    -- The example design uses Block RAM based frame generators to provide test
    -- data to the GTXs for transmission. By default the frame generators are 
    -- loaded with an incrementing data sequence that includes commas/alignment
    -- characters for alignment. If your protocol uses channel bonding, the 
    -- frame generator will also be preloaded with a channel bonding sequence.
    
    -- You can modify the data transmitted by changing the INIT values of the frame
    -- generator in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.

    tile0_frame_gen0 : FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        MEM_00                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_01                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_02                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_03                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_04                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_05                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_06                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_07                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_08                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_09                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_0A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_0B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_0C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_0D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_0E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_0F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_10                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_11                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_12                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_13                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_14                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_15                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_16                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_17                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_18                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_19                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_1A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_1B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_1C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_1D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_1E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_1F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_20                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_21                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_22                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_23                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_24                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_25                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_26                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_27                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_28                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_29                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_2A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_2B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_2C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_2D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_2E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_2F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_30                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_31                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_32                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_33                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_34                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_35                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_36                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_37                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_38                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_39                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_3A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_3B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_3C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_3D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_3E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_3F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000010"
    )
    port map
    (
        -- User Interface
        TX_DATA(39 downto 20)           =>      tile0_txdata0_float_i,
        TX_DATA(19 downto 0)            =>      tile0_txdata0_i,
        TX_CHARISK                      =>      open,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk0_i,
        SYSTEM_RESET                    =>      tile0_tx_system_reset0_c
    );
    
    tile0_frame_gen1 : FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        MEM_00                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_01                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_02                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_03                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_04                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_05                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_06                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_07                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_08                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_09                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_0A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_0B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_0C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_0D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_0E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_0F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_10                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_11                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_12                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_13                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_14                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_15                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_16                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_17                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_18                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_19                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_1A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_1B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_1C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_1D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_1E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_1F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_20                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_21                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_22                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_23                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_24                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_25                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_26                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_27                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_28                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_29                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_2A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_2B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_2C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_2D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_2E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_2F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_30                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_31                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_32                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_33                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_34                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_35                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_36                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_37                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_38                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_39                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_3A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_3B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_3C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_3D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_3E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_3F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000010"
    )
    port map
    (
        -- User Interface
        TX_DATA(39 downto 20)           =>      tile0_txdata1_float_i,
        TX_DATA(19 downto 0)            =>      tile0_txdata1_i,
        TX_CHARISK                      =>      open,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk0_i,
        SYSTEM_RESET                    =>      tile0_tx_system_reset1_c
    );
    
    tile1_frame_gen0 : FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        MEM_00                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_01                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_02                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_03                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_04                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_05                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_06                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_07                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_08                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_09                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_0A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_0B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_0C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_0D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_0E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_0F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_10                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_11                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_12                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_13                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_14                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_15                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_16                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_17                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_18                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_19                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_1A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_1B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_1C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_1D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_1E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_1F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_20                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_21                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_22                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_23                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_24                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_25                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_26                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_27                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_28                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_29                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_2A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_2B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_2C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_2D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_2E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_2F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_30                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_31                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_32                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_33                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_34                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_35                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_36                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_37                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_38                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_39                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_3A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_3B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_3C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_3D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_3E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_3F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000010"
    )
    port map
    (
        -- User Interface
        TX_DATA(39 downto 20)           =>      tile1_txdata0_float_i,
        TX_DATA(19 downto 0)            =>      tile1_txdata0_i,
        TX_CHARISK                      =>      open,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk0_i,
        SYSTEM_RESET                    =>      tile1_tx_system_reset0_c
    );
    
    tile1_frame_gen1 : FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        MEM_00                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_01                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_02                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_03                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_04                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_05                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_06                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_07                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_08                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_09                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_0A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_0B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_0C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_0D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_0E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_0F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_10                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_11                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_12                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_13                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_14                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_15                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_16                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_17                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_18                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_19                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_1A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_1B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_1C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_1D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_1E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_1F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_20                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_21                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_22                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_23                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_24                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_25                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_26                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_27                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_28                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_29                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_2A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_2B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_2C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_2D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_2E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_2F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_30                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_31                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_32                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_33                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_34                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_35                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_36                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_37                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_38                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_39                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_3A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_3B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_3C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_3D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_3E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_3F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000010"
    )
    port map
    (
        -- User Interface
        TX_DATA(39 downto 20)           =>      tile1_txdata1_float_i,
        TX_DATA(19 downto 0)            =>      tile1_txdata1_i,
        TX_CHARISK                      =>      open,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk0_i,
        SYSTEM_RESET                    =>      tile1_tx_system_reset1_c
    );
    
    tile2_frame_gen0 : FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        MEM_00                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_01                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_02                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_03                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_04                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_05                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_06                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_07                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_08                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_09                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_0A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_0B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_0C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_0D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_0E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_0F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_10                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_11                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_12                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_13                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_14                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_15                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_16                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_17                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_18                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_19                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_1A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_1B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_1C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_1D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_1E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_1F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_20                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_21                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_22                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_23                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_24                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_25                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_26                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_27                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_28                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_29                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_2A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_2B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_2C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_2D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_2E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_2F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_30                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_31                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_32                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_33                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_34                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_35                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_36                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_37                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_38                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_39                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_3A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_3B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_3C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_3D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_3E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_3F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000010"
    )
    port map
    (
        -- User Interface
        TX_DATA(39 downto 20)           =>      tile2_txdata0_float_i,
        TX_DATA(19 downto 0)            =>      tile2_txdata0_i,
        TX_CHARISK                      =>      open,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk0_i,
        SYSTEM_RESET                    =>      tile2_tx_system_reset0_c
    );
    
    tile2_frame_gen1 : FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        MEM_00                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_01                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_02                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_03                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_04                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_05                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_06                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_07                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_08                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_09                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_0A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_0B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_0C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_0D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_0E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_0F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_10                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_11                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_12                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_13                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_14                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_15                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_16                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_17                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_18                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_19                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_1A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_1B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_1C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_1D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_1E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_1F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_20                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_21                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_22                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_23                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_24                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_25                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_26                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_27                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_28                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_29                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_2A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_2B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_2C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_2D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_2E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_2F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_30                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_31                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_32                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_33                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_34                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_35                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_36                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_37                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEM_38                  =>  x"0000380d0000300b00002809000020070000180500001003000002bc00000400",
        MEM_39                  =>  x"0000781d0000701b00006819000060170000581500005013000048110000400f",
        MEM_3A                  =>  x"0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f",
        MEM_3B                  =>  x"0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f",
        MEM_3C                  =>  x"0001384d0001304b00012849000120470001184500011043000108410001003f",
        MEM_3D                  =>  x"0001785d0001705b00016859000160570001585500015053000148510001404f",
        MEM_3E                  =>  x"0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f",
        MEM_3F                  =>  x"0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000010"
    )
    port map
    (
        -- User Interface
        TX_DATA(39 downto 20)           =>      tile2_txdata1_float_i,
        TX_DATA(19 downto 0)            =>      tile2_txdata1_i,
        TX_CHARISK                      =>      open,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk0_i,
        SYSTEM_RESET                    =>      tile2_tx_system_reset1_c
    );
    


    ---------------------------------- Frame Checkers -------------------------
    -- The example design uses Block RAM based frame checkers to verify incoming  
    -- data. By default the frame generators are loaded with a data sequence that 
    -- matches the outgoing sequence of the frame generators for the TX ports.
    
    -- You can modify the expected data sequence by changing the INIT values of the frame
    -- checkers in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.
    
    -- When the frame checker receives data, it attempts to synchronise to the 
    -- incoming pattern by looking for the first sequence in the pattern. Once it 
    -- finds the first sequence, it increments through the sequence, and indicates an 
    -- error whenever the next value received does not match the expected value.

    tile0_frame_check0_reset_i              <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else tile0_matchn0_i;

    -- tile0_frame_check0 is always connected to the lane with the start of char
    -- and this lane starts off the data checking on all the other lanes. The INC_IN port is tied off
    tile0_inc_in0_i                         <= '0';

    tile0_frame_check0 : FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      16,
        USE_COMMA                       =>      1,
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        CONFIG_INDEPENDENT_LANES        =>      1,
        START_OF_PACKET_CHAR            =>      x"bc",
        MEM_00                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_01                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_02                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_03                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_04                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_05                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_06                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_07                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_08                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_09                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_0A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_0B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_0C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_0D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_0E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_0F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_10                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_11                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_12                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_13                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_14                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_15                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_16                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_17                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_18                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_19                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_1A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_1B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_1C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_1D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_1E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_1F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_20                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_21                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_22                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_23                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_24                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_25                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_26                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_27                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_28                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_29                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_2A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_2B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_2C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_2D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_2E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_2F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_30                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_31                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_32                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_33                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_34                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_35                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_36                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_37                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_38                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_39                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_3A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_3B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_3C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_3D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_3E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_3F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000010"
    )
    port map
    (
        -- MGT Interface
        RX_DATA                         =>      tile0_rxdata0_i,
        RX_ENMCOMMA_ALIGN               =>      tile0_rxenmcommaalign0_i,
        RX_ENPCOMMA_ALIGN               =>      tile0_rxenpcommaalign0_i,
        RX_ENCHAN_SYNC                  =>      open,
        RX_CHANBOND_SEQ                 =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      tile0_inc_in0_i,
        INC_OUT                         =>      tile0_inc_out0_i,
        PATTERN_MATCH_N                 =>      tile0_matchn0_i,
        RESET_ON_ERROR                  =>      tile0_frame_check0_reset_i,
        -- System Interface
        USER_CLK                        =>      tile0_rxusrclk0_i,
        SYSTEM_RESET                    =>      tile0_rx_system_reset0_c,
        ERROR_COUNT                     =>      tile0_error_count0_i
    );
        
    tile0_frame_check1_reset_i              <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else tile0_matchn1_i;

    -- tile0_frame_check0 is always connected to the lane with the start of char
    -- and this lane starts off the data checking on all the other lanes. The INC_IN port is tied off
    tile0_inc_in1_i                         <= '0';

    tile0_frame_check1 : FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      16,
        USE_COMMA                       =>      1,
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        CONFIG_INDEPENDENT_LANES        =>      1,
        START_OF_PACKET_CHAR            =>      x"bc",
        MEM_00                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_01                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_02                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_03                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_04                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_05                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_06                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_07                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_08                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_09                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_0A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_0B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_0C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_0D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_0E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_0F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_10                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_11                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_12                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_13                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_14                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_15                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_16                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_17                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_18                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_19                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_1A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_1B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_1C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_1D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_1E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_1F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_20                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_21                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_22                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_23                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_24                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_25                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_26                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_27                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_28                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_29                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_2A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_2B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_2C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_2D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_2E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_2F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_30                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_31                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_32                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_33                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_34                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_35                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_36                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_37                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_38                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_39                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_3A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_3B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_3C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_3D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_3E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_3F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000010"
    )
    port map
    (
        -- MGT Interface
        RX_DATA                         =>      tile0_rxdata1_i,
        RX_ENMCOMMA_ALIGN               =>      tile0_rxenmcommaalign1_i,
        RX_ENPCOMMA_ALIGN               =>      tile0_rxenpcommaalign1_i,
        RX_ENCHAN_SYNC                  =>      open,
        RX_CHANBOND_SEQ                 =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      tile0_inc_in1_i,
        INC_OUT                         =>      tile0_inc_out1_i,
        PATTERN_MATCH_N                 =>      tile0_matchn1_i,
        RESET_ON_ERROR                  =>      tile0_frame_check1_reset_i,
        -- System Interface
        USER_CLK                        =>      tile0_rxusrclk1_i,
        SYSTEM_RESET                    =>      tile0_rx_system_reset1_c,
        ERROR_COUNT                     =>      tile0_error_count1_i
    );
        
    tile1_frame_check0_reset_i              <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else tile1_matchn0_i;

    -- in the "independent lanes" configuration, each of the lanes looks for the unique start char and
    -- in this case, the INC_IN port is tied off.
    -- Else, the data checking is triggered by the "master" lane
    tile1_inc_in0_i                         <= tile0_inc_out0_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else '0';

    tile1_frame_check0 : FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      16,
        USE_COMMA                       =>      1,
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        CONFIG_INDEPENDENT_LANES        =>      EXAMPLE_CONFIG_INDEPENDENT_LANES,
        START_OF_PACKET_CHAR            =>      x"bc",
        MEM_00                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_01                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_02                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_03                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_04                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_05                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_06                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_07                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_08                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_09                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_0A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_0B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_0C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_0D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_0E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_0F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_10                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_11                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_12                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_13                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_14                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_15                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_16                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_17                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_18                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_19                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_1A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_1B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_1C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_1D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_1E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_1F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_20                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_21                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_22                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_23                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_24                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_25                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_26                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_27                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_28                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_29                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_2A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_2B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_2C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_2D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_2E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_2F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_30                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_31                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_32                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_33                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_34                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_35                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_36                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_37                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_38                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_39                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_3A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_3B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_3C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_3D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_3E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_3F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000010"
    )
    port map
    (
        -- MGT Interface
        RX_DATA                         =>      tile1_rxdata0_i,
        RX_ENMCOMMA_ALIGN               =>      tile1_rxenmcommaalign0_i,
        RX_ENPCOMMA_ALIGN               =>      tile1_rxenpcommaalign0_i,
        RX_ENCHAN_SYNC                  =>      open,
        RX_CHANBOND_SEQ                 =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      tile1_inc_in0_i,
        INC_OUT                         =>      tile1_inc_out0_i,
        PATTERN_MATCH_N                 =>      tile1_matchn0_i,
        RESET_ON_ERROR                  =>      tile1_frame_check0_reset_i,
        -- System Interface
        USER_CLK                        =>      tile1_rxusrclk0_i,
        SYSTEM_RESET                    =>      tile1_rx_system_reset0_c,
        ERROR_COUNT                     =>      tile1_error_count0_i
    );
        
    tile1_frame_check1_reset_i              <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else tile1_matchn1_i;

    -- in the "independent lanes" configuration, each of the lanes looks for the unique start char and
    -- in this case, the INC_IN port is tied off.
    -- Else, the data checking is triggered by the "master" lane
    tile1_inc_in1_i                         <= tile0_inc_out1_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else '0';

    tile1_frame_check1 : FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      16,
        USE_COMMA                       =>      1,
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        CONFIG_INDEPENDENT_LANES        =>      EXAMPLE_CONFIG_INDEPENDENT_LANES,
        START_OF_PACKET_CHAR            =>      x"bc",
        MEM_00                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_01                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_02                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_03                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_04                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_05                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_06                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_07                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_08                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_09                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_0A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_0B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_0C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_0D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_0E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_0F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_10                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_11                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_12                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_13                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_14                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_15                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_16                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_17                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_18                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_19                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_1A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_1B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_1C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_1D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_1E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_1F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_20                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_21                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_22                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_23                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_24                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_25                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_26                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_27                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_28                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_29                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_2A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_2B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_2C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_2D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_2E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_2F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_30                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_31                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_32                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_33                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_34                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_35                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_36                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_37                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_38                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_39                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_3A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_3B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_3C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_3D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_3E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_3F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000010"
    )
    port map
    (
        -- MGT Interface
        RX_DATA                         =>      tile1_rxdata1_i,
        RX_ENMCOMMA_ALIGN               =>      tile1_rxenmcommaalign1_i,
        RX_ENPCOMMA_ALIGN               =>      tile1_rxenpcommaalign1_i,
        RX_ENCHAN_SYNC                  =>      open,
        RX_CHANBOND_SEQ                 =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      tile1_inc_in1_i,
        INC_OUT                         =>      tile1_inc_out1_i,
        PATTERN_MATCH_N                 =>      tile1_matchn1_i,
        RESET_ON_ERROR                  =>      tile1_frame_check1_reset_i,
        -- System Interface
        USER_CLK                        =>      tile1_rxusrclk1_i,
        SYSTEM_RESET                    =>      tile1_rx_system_reset1_c,
        ERROR_COUNT                     =>      tile1_error_count1_i
    );
        
    tile2_frame_check0_reset_i              <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else tile2_matchn0_i;

    -- in the "independent lanes" configuration, each of the lanes looks for the unique start char and
    -- in this case, the INC_IN port is tied off.
    -- Else, the data checking is triggered by the "master" lane
    tile2_inc_in0_i                         <= tile0_inc_out0_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else '0';

    tile2_frame_check0 : FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      16,
        USE_COMMA                       =>      1,
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        CONFIG_INDEPENDENT_LANES        =>      EXAMPLE_CONFIG_INDEPENDENT_LANES,
        START_OF_PACKET_CHAR            =>      x"bc",
        MEM_00                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_01                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_02                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_03                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_04                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_05                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_06                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_07                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_08                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_09                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_0A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_0B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_0C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_0D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_0E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_0F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_10                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_11                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_12                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_13                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_14                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_15                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_16                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_17                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_18                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_19                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_1A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_1B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_1C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_1D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_1E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_1F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_20                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_21                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_22                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_23                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_24                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_25                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_26                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_27                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_28                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_29                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_2A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_2B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_2C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_2D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_2E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_2F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_30                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_31                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_32                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_33                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_34                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_35                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_36                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_37                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_38                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_39                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_3A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_3B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_3C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_3D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_3E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_3F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000010"
    )
    port map
    (
        -- MGT Interface
        RX_DATA                         =>      tile2_rxdata0_i,
        RX_ENMCOMMA_ALIGN               =>      tile2_rxenmcommaalign0_i,
        RX_ENPCOMMA_ALIGN               =>      tile2_rxenpcommaalign0_i,
        RX_ENCHAN_SYNC                  =>      open,
        RX_CHANBOND_SEQ                 =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      tile2_inc_in0_i,
        INC_OUT                         =>      tile2_inc_out0_i,
        PATTERN_MATCH_N                 =>      tile2_matchn0_i,
        RESET_ON_ERROR                  =>      tile2_frame_check0_reset_i,
        -- System Interface
        USER_CLK                        =>      tile2_rxusrclk0_i,
        SYSTEM_RESET                    =>      tile2_rx_system_reset0_c,
        ERROR_COUNT                     =>      tile2_error_count0_i
    );
        
    tile2_frame_check1_reset_i              <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else tile2_matchn1_i;

    -- in the "independent lanes" configuration, each of the lanes looks for the unique start char and
    -- in this case, the INC_IN port is tied off.
    -- Else, the data checking is triggered by the "master" lane
    tile2_inc_in1_i                         <= tile0_inc_out1_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else '0';

    tile2_frame_check1 : FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      16,
        USE_COMMA                       =>      1,
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        CONFIG_INDEPENDENT_LANES        =>      EXAMPLE_CONFIG_INDEPENDENT_LANES,
        START_OF_PACKET_CHAR            =>      x"bc",
        MEM_00                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_01                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_02                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_03                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_04                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_05                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_06                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_07                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_08                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_09                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_0A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_0B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_0C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_0D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_0E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_0F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_10                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_11                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_12                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_13                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_14                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_15                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_16                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_17                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_18                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_19                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_1A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_1B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_1C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_1D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_1E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_1F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_20                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_21                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_22                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_23                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_24                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_25                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_26                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_27                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_28                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_29                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_2A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_2B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_2C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_2D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_2E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_2F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_30                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_31                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_32                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_33                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_34                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_35                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_36                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_37                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEM_38                  =>  x"00000e0d00000c0b00000a09000008070000060500000403000002bc00000100",
        MEM_39                  =>  x"00001e1d00001c1b00001a19000018170000161500001413000012110000100f",
        MEM_3A                  =>  x"00002e2d00002c2b00002a29000028270000262500002423000022210000201f",
        MEM_3B                  =>  x"00003e3d00003c3b00003a39000038370000363500003433000032310000302f",
        MEM_3C                  =>  x"00004e4d00004c4b00004a49000048470000464500004443000042410000403f",
        MEM_3D                  =>  x"00005e5d00005c5b00005a59000058570000565500005453000052510000504f",
        MEM_3E                  =>  x"00006e6d00006c6b00006a69000068670000666500006463000062610000605f",
        MEM_3F                  =>  x"00007e7d00007c7b00007a79000078770000767500007473000072710000706f",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000010",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000010"
    )
    port map
    (
        -- MGT Interface
        RX_DATA                         =>      tile2_rxdata1_i,
        RX_ENMCOMMA_ALIGN               =>      tile2_rxenmcommaalign1_i,
        RX_ENPCOMMA_ALIGN               =>      tile2_rxenpcommaalign1_i,
        RX_ENCHAN_SYNC                  =>      open,
        RX_CHANBOND_SEQ                 =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      tile2_inc_in1_i,
        INC_OUT                         =>      tile2_inc_out1_i,
        PATTERN_MATCH_N                 =>      tile2_matchn1_i,
        RESET_ON_ERROR                  =>      tile2_frame_check1_reset_i,
        -- System Interface
        USER_CLK                        =>      tile2_rxusrclk1_i,
        SYSTEM_RESET                    =>      tile2_rx_system_reset1_c,
        ERROR_COUNT                     =>      tile2_error_count1_i
    );
        





    ----------------------------- Chipscope Connections -----------------------
    -- When the example design is run in hardware, it uses chipscope to allow the
    -- example design and GTX wrapper to be controlled and monitored. The 
    -- EXAMPLE_USE_CHIPSCOPE parameter allows chipscope to be removed for simulation.
    
chipscope : if EXAMPLE_USE_CHIPSCOPE = 1 generate


    -- Shared VIO for all tiles
    shared_vio_i : shared_vio
    port map
    (
        control                         =>      shared_vio_control_i,
        async_in                        =>      shared_vio_in_i,
        async_out                       =>      shared_vio_out_i
    );

    -- ICON for all VIOs 
    i_icon : icon
    port map
    (
        control0                        =>      shared_vio_control_i,
        control1                        =>      tx_data_vio_control0_i,
        control2                        =>      rx_data_vio_control0_i,
        control3                        =>      ila_control0_i,
        control4                        =>      tx_data_vio_control1_i,
        control5                        =>      rx_data_vio_control1_i,
        control6                        =>      ila_control1_i
    );

    -- TX VIO 
    tx_data_vio0_i : shared_vio
    port map
    (
        control                         =>      tx_data_vio_control0_i,
        async_in                        =>      tx_data_vio_in0_i,
        async_out                       =>      tx_data_vio_out0_i
    );
    
    -- RX VIO 
    rx_data_vio0_i : shared_vio
    port map
    (
        control                         =>      rx_data_vio_control0_i,
        async_in                        =>      rx_data_vio_in0_i,
        async_out                       =>      rx_data_vio_out0_i
    );
    
    -- RX ILA
    ila0_i : ila
    port map
    (
        control                         =>      ila_control0_i,
        clk                             =>      ila_clk0_i,
        trig0                           =>      ila_in0_i
    );

    
    -- The RX ILA must use the same clock as the selected transceiver
    process(mux_sel_i)
    begin
      case mux_sel_i is
        when "00" => async_mux0_sel_i <= "00";
        when "01" => async_mux0_sel_i <= "01";
        when "10" => async_mux0_sel_i <= "10";
        when others => async_mux0_sel_i <= "00";
      end case;
    end process;

    not_async_mux0_sel_i <= not async_mux0_sel_i;

    async_mux0_inst0: BUFGCTRL
    port map
    (
        O => ila_clk0_mux_out0_i,
        I0 => tile0_rxusrclk0_i,
        I1 => tile1_rxusrclk0_i,
        CE0 => '1',
        CE1 => '1',
        S0 => not_async_mux0_sel_i(0),
        S1 => async_mux0_sel_i(0),
        IGNORE0 => '1',
        IGNORE1 => '1'
    );

    async_mux0_inst1: BUFGCTRL
    port map
    (
        O => ila_clk0_i,
        I0 => ila_clk0_mux_out0_i,
        I1 => tile2_rxusrclk0_i,
        CE0 => '1',
        CE1 => '1',
        S0 => not_async_mux0_sel_i(1),
        S1 => async_mux0_sel_i(1),
        IGNORE0 => '1',
        IGNORE1 => '1'
    );



    -- TX VIO 
    tx_data_vio1_i : shared_vio
    port map
    (
        control                         =>      tx_data_vio_control1_i,
        async_in                        =>      tx_data_vio_in1_i,
        async_out                       =>      tx_data_vio_out1_i
    );
    
    -- RX VIO 
    rx_data_vio1_i : shared_vio
    port map
    (
        control                         =>      rx_data_vio_control1_i,
        async_in                        =>      rx_data_vio_in1_i,
        async_out                       =>      rx_data_vio_out1_i
    );
    
    -- RX ILA
    ila1_i : ila
    port map
    (
        control                         =>      ila_control1_i,
        clk                             =>      ila_clk1_i,
        trig0                           =>      ila_in1_i
    );

    
    -- The RX ILA must use the same clock as the selected transceiver
    process(mux_sel_i)
    begin
      case mux_sel_i is
        when "00" => async_mux1_sel_i <= "00";
        when "01" => async_mux1_sel_i <= "01";
        when "10" => async_mux1_sel_i <= "10";
        when others => async_mux1_sel_i <= "00";
      end case;
    end process;

    not_async_mux1_sel_i <= not async_mux1_sel_i;

    async_mux1_inst0: BUFGCTRL
    port map
    (
        O => ila_clk1_mux_out0_i,
        I0 => tile0_rxusrclk1_i,
        I1 => tile1_rxusrclk1_i,
        CE0 => '1',
        CE1 => '1',
        S0 => not_async_mux1_sel_i(0),
        S1 => async_mux1_sel_i(0),
        IGNORE0 => '1',
        IGNORE1 => '1'
    );

    async_mux1_inst1: BUFGCTRL
    port map
    (
        O => ila_clk1_i,
        I0 => ila_clk1_mux_out0_i,
        I1 => tile2_rxusrclk1_i,
        CE0 => '1',
        CE1 => '1',
        S0 => not_async_mux1_sel_i(1),
        S1 => async_mux1_sel_i(1),
        IGNORE0 => '1',
        IGNORE1 => '1'
    );




    -- assign resets for frame_gen modules
    tile0_tx_system_reset0_c                <= not tile0_tx_resetdone0_r2 or user_tx_reset_i;
    tile0_tx_system_reset1_c                <= not tile0_tx_resetdone1_r2 or user_tx_reset_i;
    tile1_tx_system_reset0_c                <= not tile1_tx_resetdone0_r2 or user_tx_reset_i;
    tile1_tx_system_reset1_c                <= not tile1_tx_resetdone1_r2 or user_tx_reset_i;
    tile2_tx_system_reset0_c                <= not tile2_tx_resetdone0_r2 or user_tx_reset_i;
    tile2_tx_system_reset1_c                <= not tile2_tx_resetdone1_r2 or user_tx_reset_i;
    -- assign resets for frame_check modules
    tile0_rx_system_reset0_c                <= not tile0_rx_resetdone0_r2 or user_rx_reset_i;
    tile0_rx_system_reset1_c                <= not tile0_rx_resetdone1_r2 or user_rx_reset_i;
    tile1_rx_system_reset0_c                <= not tile1_rx_resetdone0_r2 or user_rx_reset_i;
    tile1_rx_system_reset1_c                <= not tile1_rx_resetdone1_r2 or user_rx_reset_i;
    tile2_rx_system_reset0_c                <= not tile2_rx_resetdone0_r2 or user_rx_reset_i;
    tile2_rx_system_reset1_c                <= not tile2_rx_resetdone1_r2 or user_rx_reset_i;


    tile0_gtxreset_i                        <= gtxreset_i;
    tile1_gtxreset_i                        <= gtxreset_i;
    tile2_gtxreset_i                        <= gtxreset_i;

    -- Shared VIO Outputs
    gtxreset_i                              <= shared_vio_out_i(31);
    user_tx_reset_i                         <= shared_vio_out_i(30);
    user_rx_reset_i                         <= shared_vio_out_i(29);
    mux_sel_i                               <= shared_vio_out_i(28 downto 27);

    -- Shared VIO Inputs
    shared_vio_in_i(31)                     <= tile0_plllkdet_i;
    shared_vio_in_i(30)                     <= tile1_plllkdet_i;
    shared_vio_in_i(29)                     <= tile2_plllkdet_i;
    shared_vio_in_i(28 downto 0)            <= "00000000000000000000000000000";

    -- Chipscope connections for GTP0 on Tile 0
    tile0_tx_data_vio_in0_i(31 downto 0)    <= "00000000000000000000000000000000";
    tile0_rx_data_vio_in0_i(31)             <= tile0_resetdone0_i;
    tile0_rx_data_vio_in0_i(30 downto 0)    <= "0000000000000000000000000000000";
    tile0_rxeqmix0_i                        <= rx_data_vio_out0_i(31 downto 30);
    tile0_rxpolarity0_i                     <= rx_data_vio_out0_i(29);
    tile0_ila_in0_i(84 downto 83)           <= tile0_rxchariscomma0_i;
    tile0_ila_in0_i(82 downto 81)           <= tile0_rxdisperr0_i;
    tile0_ila_in0_i(80 downto 79)           <= tile0_rxnotintable0_i;
    tile0_ila_in0_i(78)                     <= tile0_rxbyteisaligned0_i;
    tile0_ila_in0_i(77 downto 62)           <= tile0_rxdata0_i;
    tile0_ila_in0_i(61 downto 54)           <= tile0_error_count0_i;
    tile0_ila_in0_i(53 downto 0)            <= "000000000000000000000000000000000000000000000000000000";

    -- Chipscope connections for GTP1 on Tile 0
    tile0_tx_data_vio_in1_i(31 downto 0)    <= "00000000000000000000000000000000";
    tile0_rx_data_vio_in1_i(31)             <= tile0_resetdone1_i;
    tile0_rx_data_vio_in1_i(30 downto 0)    <= "0000000000000000000000000000000";
    tile0_rxeqmix1_i                        <= rx_data_vio_out1_i(31 downto 30);
    tile0_rxpolarity1_i                     <= rx_data_vio_out1_i(29);
    tile0_ila_in1_i(84 downto 83)           <= tile0_rxchariscomma1_i;
    tile0_ila_in1_i(82 downto 81)           <= tile0_rxdisperr1_i;
    tile0_ila_in1_i(80 downto 79)           <= tile0_rxnotintable1_i;
    tile0_ila_in1_i(78)                     <= tile0_rxbyteisaligned1_i;
    tile0_ila_in1_i(77 downto 62)           <= tile0_rxdata1_i;
    tile0_ila_in1_i(61 downto 54)           <= tile0_error_count1_i;
    tile0_ila_in1_i(53 downto 0)            <= "000000000000000000000000000000000000000000000000000000";

    -- Chipscope connections for GTP0 on Tile 1
    tile1_tx_data_vio_in0_i(31 downto 0)    <= "00000000000000000000000000000000";
    tile1_rx_data_vio_in0_i(31)             <= tile1_resetdone0_i;
    tile1_rx_data_vio_in0_i(30 downto 0)    <= "0000000000000000000000000000000";
    tile1_rxeqmix0_i                        <= rx_data_vio_out0_i(31 downto 30);
    tile1_rxpolarity0_i                     <= rx_data_vio_out0_i(29);
    tile1_ila_in0_i(84 downto 83)           <= tile1_rxchariscomma0_i;
    tile1_ila_in0_i(82 downto 81)           <= tile1_rxdisperr0_i;
    tile1_ila_in0_i(80 downto 79)           <= tile1_rxnotintable0_i;
    tile1_ila_in0_i(78)                     <= tile1_rxbyteisaligned0_i;
    tile1_ila_in0_i(77 downto 62)           <= tile1_rxdata0_i;
    tile1_ila_in0_i(61 downto 54)           <= tile1_error_count0_i;
    tile1_ila_in0_i(53 downto 0)            <= "000000000000000000000000000000000000000000000000000000";

    -- Chipscope connections for GTP1 on Tile 1
    tile1_tx_data_vio_in1_i(31 downto 0)    <= "00000000000000000000000000000000";
    tile1_rx_data_vio_in1_i(31)             <= tile1_resetdone1_i;
    tile1_rx_data_vio_in1_i(30 downto 0)    <= "0000000000000000000000000000000";
    tile1_rxeqmix1_i                        <= rx_data_vio_out1_i(31 downto 30);
    tile1_rxpolarity1_i                     <= rx_data_vio_out1_i(29);
    tile1_ila_in1_i(84 downto 83)           <= tile1_rxchariscomma1_i;
    tile1_ila_in1_i(82 downto 81)           <= tile1_rxdisperr1_i;
    tile1_ila_in1_i(80 downto 79)           <= tile1_rxnotintable1_i;
    tile1_ila_in1_i(78)                     <= tile1_rxbyteisaligned1_i;
    tile1_ila_in1_i(77 downto 62)           <= tile1_rxdata1_i;
    tile1_ila_in1_i(61 downto 54)           <= tile1_error_count1_i;
    tile1_ila_in1_i(53 downto 0)            <= "000000000000000000000000000000000000000000000000000000";

    -- Chipscope connections for GTP0 on Tile 2
    tile2_tx_data_vio_in0_i(31 downto 0)    <= "00000000000000000000000000000000";
    tile2_rx_data_vio_in0_i(31)             <= tile2_resetdone0_i;
    tile2_rx_data_vio_in0_i(30 downto 0)    <= "0000000000000000000000000000000";
    tile2_rxeqmix0_i                        <= rx_data_vio_out0_i(31 downto 30);
    tile2_rxpolarity0_i                     <= rx_data_vio_out0_i(29);
    tile2_ila_in0_i(84 downto 83)           <= tile2_rxchariscomma0_i;
    tile2_ila_in0_i(82 downto 81)           <= tile2_rxdisperr0_i;
    tile2_ila_in0_i(80 downto 79)           <= tile2_rxnotintable0_i;
    tile2_ila_in0_i(78)                     <= tile2_rxbyteisaligned0_i;
    tile2_ila_in0_i(77 downto 62)           <= tile2_rxdata0_i;
    tile2_ila_in0_i(61 downto 54)           <= tile2_error_count0_i;
    tile2_ila_in0_i(53 downto 0)            <= "000000000000000000000000000000000000000000000000000000";

    -- Chipscope connections for GTP1 on Tile 2
    tile2_tx_data_vio_in1_i(31 downto 0)    <= "00000000000000000000000000000000";
    tile2_rx_data_vio_in1_i(31)             <= tile2_resetdone1_i;
    tile2_rx_data_vio_in1_i(30 downto 0)    <= "0000000000000000000000000000000";
    tile2_rxeqmix1_i                        <= rx_data_vio_out1_i(31 downto 30);
    tile2_rxpolarity1_i                     <= rx_data_vio_out1_i(29);
    tile2_ila_in1_i(84 downto 83)           <= tile2_rxchariscomma1_i;
    tile2_ila_in1_i(82 downto 81)           <= tile2_rxdisperr1_i;
    tile2_ila_in1_i(80 downto 79)           <= tile2_rxnotintable1_i;
    tile2_ila_in1_i(78)                     <= tile2_rxbyteisaligned1_i;
    tile2_ila_in1_i(77 downto 62)           <= tile2_rxdata1_i;
    tile2_ila_in1_i(61 downto 54)           <= tile2_error_count1_i;
    tile2_ila_in1_i(53 downto 0)            <= "000000000000000000000000000000000000000000000000000000";


    --Mux inputs to Chipscope modules based on mux_sel_i
    tx_data_vio_in0_i                   <=      tile0_tx_data_vio_in0_i when (mux_sel_i = "00")
                                        else    tile1_tx_data_vio_in0_i when (mux_sel_i = "01")
                                        else    tile2_tx_data_vio_in0_i;


    rx_data_vio_in0_i                   <=      tile0_rx_data_vio_in0_i when (mux_sel_i = "00")
                                        else    tile1_rx_data_vio_in0_i when (mux_sel_i = "01")
                                        else    tile2_rx_data_vio_in0_i;


    ila_in0_i                           <=      tile0_ila_in0_i when (mux_sel_i = "00")
                                        else    tile1_ila_in0_i when (mux_sel_i = "01")
                                        else    tile2_ila_in0_i;



    tx_data_vio_in1_i                   <=      tile0_tx_data_vio_in1_i when (mux_sel_i = "00")
                                        else    tile1_tx_data_vio_in1_i when (mux_sel_i = "01")
                                        else    tile2_tx_data_vio_in1_i;


    rx_data_vio_in1_i                   <=      tile0_rx_data_vio_in1_i when (mux_sel_i = "00")
                                        else    tile1_rx_data_vio_in1_i when (mux_sel_i = "01")
                                        else    tile2_rx_data_vio_in1_i;


    ila_in1_i                           <=      tile0_ila_in1_i when (mux_sel_i = "00")
                                        else    tile1_ila_in1_i when (mux_sel_i = "01")
                                        else    tile2_ila_in1_i;





   
end generate chipscope;


no_chipscope : if EXAMPLE_USE_CHIPSCOPE = 0 generate

    -- If Chipscope is not being used, drive GTX reset signal
    -- from the top level ports
    tile0_gtxreset_i                        <= GTXRESET_IN;
    tile1_gtxreset_i                        <= GTXRESET_IN;
    tile2_gtxreset_i                        <= GTXRESET_IN;

    -- assign resets for frame_gen modules
    tile0_tx_system_reset0_c                <= not tile0_tx_resetdone0_r2;
    tile0_tx_system_reset1_c                <= not tile0_tx_resetdone1_r2;
    tile1_tx_system_reset0_c                <= not tile1_tx_resetdone0_r2;
    tile1_tx_system_reset1_c                <= not tile1_tx_resetdone1_r2;
    tile2_tx_system_reset0_c                <= not tile2_tx_resetdone0_r2;
    tile2_tx_system_reset1_c                <= not tile2_tx_resetdone1_r2;
    -- assign resets for frame_check modules
    tile0_rx_system_reset0_c                <= not tile0_rx_resetdone0_r2;
    tile0_rx_system_reset1_c                <= not tile0_rx_resetdone1_r2;
    tile1_rx_system_reset0_c                <= not tile1_rx_resetdone0_r2;
    tile1_rx_system_reset1_c                <= not tile1_rx_resetdone1_r2;
    tile2_rx_system_reset0_c                <= not tile2_rx_resetdone0_r2;
    tile2_rx_system_reset1_c                <= not tile2_rx_resetdone1_r2;

    gtxreset_i                              <= tied_to_ground_i;
    user_tx_reset_i                         <= tied_to_ground_i;
    user_rx_reset_i                         <= tied_to_ground_i;
    mux_sel_i                               <= tied_to_ground_vec_i(1 downto 0);
    tile0_rxeqmix0_i                        <= tied_to_ground_vec_i(1 downto 0);
    tile0_rxpolarity0_i                     <= tied_to_ground_i;
    tile0_rxeqmix1_i                        <= tied_to_ground_vec_i(1 downto 0);
    tile0_rxpolarity1_i                     <= tied_to_ground_i;
    tile1_rxeqmix0_i                        <= tied_to_ground_vec_i(1 downto 0);
    tile1_rxpolarity0_i                     <= tied_to_ground_i;
    tile1_rxeqmix1_i                        <= tied_to_ground_vec_i(1 downto 0);
    tile1_rxpolarity1_i                     <= tied_to_ground_i;
    tile2_rxeqmix0_i                        <= tied_to_ground_vec_i(1 downto 0);
    tile2_rxpolarity0_i                     <= tied_to_ground_i;
    tile2_rxeqmix1_i                        <= tied_to_ground_vec_i(1 downto 0);
    tile2_rxpolarity1_i                     <= tied_to_ground_i;



end generate no_chipscope;


end RTL;


