//////////////////////////////////////////////////////////////////////////////
//$Date: 2008/05/30 00:57:53 $
//$RCSfile: multi_mgt_wrapper.ejava,v $
//$Revision: 1.1.2.1 $
///////////////////////////////////////////////////////////////////////////////
//   ____  ____ 
//  /   /\/   / 
// /___/  \  /    Vendor: Xilinx 
// \   \   \/     Version : 1.5 
//  \   \         Application : RocketIO GTX Wizard 
//  /   /         Filename : gtx.v
// /___/   /\     Timestamp : 02/08/2005 09:12:43
// \   \  /  \ 
//  \___\/\___\ 
//
//
// Module GTX (a GTX Wrapper)
// Generated by Xilinx RocketIO GTX Wizard



`timescale 1ns / 1ps


//***************************** Entity Declaration ****************************

module GTX #
(
    // Simulation attributes
    parameter   WRAPPER_SIM_MODE                = "FAST",   // Set to Fast Functional Simulation Model
    parameter   WRAPPER_SIM_GTXRESET_SPEEDUP    = 0,    // Set to 1 to speed up sim reset
    parameter   WRAPPER_SIM_PLL_PERDIV2         = 9'h0fa   // Set to the VCO Unit Interval time    
)
(
    
    //_________________________________________________________________________
    //_________________________________________________________________________
    //TILE0  (Location)

    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    TILE0_RXCHARISCOMMA0_OUT,
    TILE0_RXCHARISCOMMA1_OUT,
    TILE0_RXDISPERR0_OUT,
    TILE0_RXDISPERR1_OUT,
    TILE0_RXNOTINTABLE0_OUT,
    TILE0_RXNOTINTABLE1_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    TILE0_RXBYTEISALIGNED0_OUT,
    TILE0_RXBYTEISALIGNED1_OUT,
    TILE0_RXENMCOMMAALIGN0_IN,
    TILE0_RXENMCOMMAALIGN1_IN,
    TILE0_RXENPCOMMAALIGN0_IN,
    TILE0_RXENPCOMMAALIGN1_IN,
    //----------------- Receive Ports - RX Data Path interface -----------------
    TILE0_RXDATA0_OUT,
    TILE0_RXDATA1_OUT,
    TILE0_RXRECCLK0_OUT,
    TILE0_RXRECCLK1_OUT,
    TILE0_RXUSRCLK0_IN,
    TILE0_RXUSRCLK1_IN,
    TILE0_RXUSRCLK20_IN,
    TILE0_RXUSRCLK21_IN,
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    TILE0_RXEQMIX0_IN,
    TILE0_RXEQMIX1_IN,
    TILE0_RXN0_IN,
    TILE0_RXN1_IN,
    TILE0_RXP0_IN,
    TILE0_RXP1_IN,
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    TILE0_RXPOLARITY0_IN,
    TILE0_RXPOLARITY1_IN,
    //------------------- Shared Ports - Tile and PLL Ports --------------------
    TILE0_CLKIN_IN,
    TILE0_GTXRESET_IN,
    TILE0_PLLLKDET_OUT,
    TILE0_REFCLKOUT_OUT,
    TILE0_RESETDONE0_OUT,
    TILE0_RESETDONE1_OUT,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    TILE0_TXDATA0_IN,
    TILE0_TXDATA1_IN,
    TILE0_TXUSRCLK0_IN,
    TILE0_TXUSRCLK1_IN,
    TILE0_TXUSRCLK20_IN,
    TILE0_TXUSRCLK21_IN,
    //------------- Transmit Ports - TX Driver and OOB signalling --------------
    TILE0_TXN0_OUT,
    TILE0_TXN1_OUT,
    TILE0_TXP0_OUT,
    TILE0_TXP1_OUT,


    
    //_________________________________________________________________________
    //_________________________________________________________________________
    //TILE1  (Location)

    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    TILE1_RXCHARISCOMMA0_OUT,
    TILE1_RXCHARISCOMMA1_OUT,
    TILE1_RXDISPERR0_OUT,
    TILE1_RXDISPERR1_OUT,
    TILE1_RXNOTINTABLE0_OUT,
    TILE1_RXNOTINTABLE1_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    TILE1_RXBYTEISALIGNED0_OUT,
    TILE1_RXBYTEISALIGNED1_OUT,
    TILE1_RXENMCOMMAALIGN0_IN,
    TILE1_RXENMCOMMAALIGN1_IN,
    TILE1_RXENPCOMMAALIGN0_IN,
    TILE1_RXENPCOMMAALIGN1_IN,
    //----------------- Receive Ports - RX Data Path interface -----------------
    TILE1_RXDATA0_OUT,
    TILE1_RXDATA1_OUT,
    TILE1_RXRECCLK0_OUT,
    TILE1_RXRECCLK1_OUT,
    TILE1_RXUSRCLK0_IN,
    TILE1_RXUSRCLK1_IN,
    TILE1_RXUSRCLK20_IN,
    TILE1_RXUSRCLK21_IN,
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    TILE1_RXEQMIX0_IN,
    TILE1_RXEQMIX1_IN,
    TILE1_RXN0_IN,
    TILE1_RXN1_IN,
    TILE1_RXP0_IN,
    TILE1_RXP1_IN,
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    TILE1_RXPOLARITY0_IN,
    TILE1_RXPOLARITY1_IN,
    //------------------- Shared Ports - Tile and PLL Ports --------------------
    TILE1_CLKIN_IN,
    TILE1_GTXRESET_IN,
    TILE1_PLLLKDET_OUT,
    TILE1_REFCLKOUT_OUT,
    TILE1_RESETDONE0_OUT,
    TILE1_RESETDONE1_OUT,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    TILE1_TXDATA0_IN,
    TILE1_TXDATA1_IN,
    TILE1_TXUSRCLK0_IN,
    TILE1_TXUSRCLK1_IN,
    TILE1_TXUSRCLK20_IN,
    TILE1_TXUSRCLK21_IN,
    //------------- Transmit Ports - TX Driver and OOB signalling --------------
    TILE1_TXN0_OUT,
    TILE1_TXN1_OUT,
    TILE1_TXP0_OUT,
    TILE1_TXP1_OUT,


    
    //_________________________________________________________________________
    //_________________________________________________________________________
    //TILE2  (Location)

    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    TILE2_RXCHARISCOMMA0_OUT,
    TILE2_RXCHARISCOMMA1_OUT,
    TILE2_RXDISPERR0_OUT,
    TILE2_RXDISPERR1_OUT,
    TILE2_RXNOTINTABLE0_OUT,
    TILE2_RXNOTINTABLE1_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    TILE2_RXBYTEISALIGNED0_OUT,
    TILE2_RXBYTEISALIGNED1_OUT,
    TILE2_RXENMCOMMAALIGN0_IN,
    TILE2_RXENMCOMMAALIGN1_IN,
    TILE2_RXENPCOMMAALIGN0_IN,
    TILE2_RXENPCOMMAALIGN1_IN,
    //----------------- Receive Ports - RX Data Path interface -----------------
    TILE2_RXDATA0_OUT,
    TILE2_RXDATA1_OUT,
    TILE2_RXRECCLK0_OUT,
    TILE2_RXRECCLK1_OUT,
    TILE2_RXUSRCLK0_IN,
    TILE2_RXUSRCLK1_IN,
    TILE2_RXUSRCLK20_IN,
    TILE2_RXUSRCLK21_IN,
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    TILE2_RXEQMIX0_IN,
    TILE2_RXEQMIX1_IN,
    TILE2_RXN0_IN,
    TILE2_RXN1_IN,
    TILE2_RXP0_IN,
    TILE2_RXP1_IN,
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    TILE2_RXPOLARITY0_IN,
    TILE2_RXPOLARITY1_IN,
    //------------------- Shared Ports - Tile and PLL Ports --------------------
    TILE2_CLKIN_IN,
    TILE2_GTXRESET_IN,
    TILE2_PLLLKDET_OUT,
    TILE2_REFCLKOUT_OUT,
    TILE2_RESETDONE0_OUT,
    TILE2_RESETDONE1_OUT,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    TILE2_TXDATA0_IN,
    TILE2_TXDATA1_IN,
    TILE2_TXUSRCLK0_IN,
    TILE2_TXUSRCLK1_IN,
    TILE2_TXUSRCLK20_IN,
    TILE2_TXUSRCLK21_IN,
    //------------- Transmit Ports - TX Driver and OOB signalling --------------
    TILE2_TXN0_OUT,
    TILE2_TXN1_OUT,
    TILE2_TXP0_OUT,
    TILE2_TXP1_OUT


);

// synthesis attribute X_CORE_INFO of GTX is "gtxwizard_v1_5, Coregen v10.1_ip3";

//***************************** Port Declarations *****************************
        


    //_________________________________________________________________________
    //_________________________________________________________________________
    //TILE0  (Location)

    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    output  [1:0]   TILE0_RXCHARISCOMMA0_OUT;
    output  [1:0]   TILE0_RXCHARISCOMMA1_OUT;
    output  [1:0]   TILE0_RXDISPERR0_OUT;
    output  [1:0]   TILE0_RXDISPERR1_OUT;
    output  [1:0]   TILE0_RXNOTINTABLE0_OUT;
    output  [1:0]   TILE0_RXNOTINTABLE1_OUT;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    output          TILE0_RXBYTEISALIGNED0_OUT;
    output          TILE0_RXBYTEISALIGNED1_OUT;
    input           TILE0_RXENMCOMMAALIGN0_IN;
    input           TILE0_RXENMCOMMAALIGN1_IN;
    input           TILE0_RXENPCOMMAALIGN0_IN;
    input           TILE0_RXENPCOMMAALIGN1_IN;
    //----------------- Receive Ports - RX Data Path interface -----------------
    output  [15:0]  TILE0_RXDATA0_OUT;
    output  [15:0]  TILE0_RXDATA1_OUT;
    output          TILE0_RXRECCLK0_OUT;
    output          TILE0_RXRECCLK1_OUT;
    input           TILE0_RXUSRCLK0_IN;
    input           TILE0_RXUSRCLK1_IN;
    input           TILE0_RXUSRCLK20_IN;
    input           TILE0_RXUSRCLK21_IN;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    input   [1:0]   TILE0_RXEQMIX0_IN;
    input   [1:0]   TILE0_RXEQMIX1_IN;
    input           TILE0_RXN0_IN;
    input           TILE0_RXN1_IN;
    input           TILE0_RXP0_IN;
    input           TILE0_RXP1_IN;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           TILE0_RXPOLARITY0_IN;
    input           TILE0_RXPOLARITY1_IN;
    //------------------- Shared Ports - Tile and PLL Ports --------------------
    input           TILE0_CLKIN_IN;
    input           TILE0_GTXRESET_IN;
    output          TILE0_PLLLKDET_OUT;
    output          TILE0_REFCLKOUT_OUT;
    output          TILE0_RESETDONE0_OUT;
    output          TILE0_RESETDONE1_OUT;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [19:0]  TILE0_TXDATA0_IN;
    input   [19:0]  TILE0_TXDATA1_IN;
    input           TILE0_TXUSRCLK0_IN;
    input           TILE0_TXUSRCLK1_IN;
    input           TILE0_TXUSRCLK20_IN;
    input           TILE0_TXUSRCLK21_IN;
    //------------- Transmit Ports - TX Driver and OOB signalling --------------
    output          TILE0_TXN0_OUT;
    output          TILE0_TXN1_OUT;
    output          TILE0_TXP0_OUT;
    output          TILE0_TXP1_OUT;



    //_________________________________________________________________________
    //_________________________________________________________________________
    //TILE1  (Location)

    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    output  [1:0]   TILE1_RXCHARISCOMMA0_OUT;
    output  [1:0]   TILE1_RXCHARISCOMMA1_OUT;
    output  [1:0]   TILE1_RXDISPERR0_OUT;
    output  [1:0]   TILE1_RXDISPERR1_OUT;
    output  [1:0]   TILE1_RXNOTINTABLE0_OUT;
    output  [1:0]   TILE1_RXNOTINTABLE1_OUT;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    output          TILE1_RXBYTEISALIGNED0_OUT;
    output          TILE1_RXBYTEISALIGNED1_OUT;
    input           TILE1_RXENMCOMMAALIGN0_IN;
    input           TILE1_RXENMCOMMAALIGN1_IN;
    input           TILE1_RXENPCOMMAALIGN0_IN;
    input           TILE1_RXENPCOMMAALIGN1_IN;
    //----------------- Receive Ports - RX Data Path interface -----------------
    output  [15:0]  TILE1_RXDATA0_OUT;
    output  [15:0]  TILE1_RXDATA1_OUT;
    output          TILE1_RXRECCLK0_OUT;
    output          TILE1_RXRECCLK1_OUT;
    input           TILE1_RXUSRCLK0_IN;
    input           TILE1_RXUSRCLK1_IN;
    input           TILE1_RXUSRCLK20_IN;
    input           TILE1_RXUSRCLK21_IN;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    input   [1:0]   TILE1_RXEQMIX0_IN;
    input   [1:0]   TILE1_RXEQMIX1_IN;
    input           TILE1_RXN0_IN;
    input           TILE1_RXN1_IN;
    input           TILE1_RXP0_IN;
    input           TILE1_RXP1_IN;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           TILE1_RXPOLARITY0_IN;
    input           TILE1_RXPOLARITY1_IN;
    //------------------- Shared Ports - Tile and PLL Ports --------------------
    input           TILE1_CLKIN_IN;
    input           TILE1_GTXRESET_IN;
    output          TILE1_PLLLKDET_OUT;
    output          TILE1_REFCLKOUT_OUT;
    output          TILE1_RESETDONE0_OUT;
    output          TILE1_RESETDONE1_OUT;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [19:0]  TILE1_TXDATA0_IN;
    input   [19:0]  TILE1_TXDATA1_IN;
    input           TILE1_TXUSRCLK0_IN;
    input           TILE1_TXUSRCLK1_IN;
    input           TILE1_TXUSRCLK20_IN;
    input           TILE1_TXUSRCLK21_IN;
    //------------- Transmit Ports - TX Driver and OOB signalling --------------
    output          TILE1_TXN0_OUT;
    output          TILE1_TXN1_OUT;
    output          TILE1_TXP0_OUT;
    output          TILE1_TXP1_OUT;



    //_________________________________________________________________________
    //_________________________________________________________________________
    //TILE2  (Location)

    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    output  [1:0]   TILE2_RXCHARISCOMMA0_OUT;
    output  [1:0]   TILE2_RXCHARISCOMMA1_OUT;
    output  [1:0]   TILE2_RXDISPERR0_OUT;
    output  [1:0]   TILE2_RXDISPERR1_OUT;
    output  [1:0]   TILE2_RXNOTINTABLE0_OUT;
    output  [1:0]   TILE2_RXNOTINTABLE1_OUT;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    output          TILE2_RXBYTEISALIGNED0_OUT;
    output          TILE2_RXBYTEISALIGNED1_OUT;
    input           TILE2_RXENMCOMMAALIGN0_IN;
    input           TILE2_RXENMCOMMAALIGN1_IN;
    input           TILE2_RXENPCOMMAALIGN0_IN;
    input           TILE2_RXENPCOMMAALIGN1_IN;
    //----------------- Receive Ports - RX Data Path interface -----------------
    output  [15:0]  TILE2_RXDATA0_OUT;
    output  [15:0]  TILE2_RXDATA1_OUT;
    output          TILE2_RXRECCLK0_OUT;
    output          TILE2_RXRECCLK1_OUT;
    input           TILE2_RXUSRCLK0_IN;
    input           TILE2_RXUSRCLK1_IN;
    input           TILE2_RXUSRCLK20_IN;
    input           TILE2_RXUSRCLK21_IN;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    input   [1:0]   TILE2_RXEQMIX0_IN;
    input   [1:0]   TILE2_RXEQMIX1_IN;
    input           TILE2_RXN0_IN;
    input           TILE2_RXN1_IN;
    input           TILE2_RXP0_IN;
    input           TILE2_RXP1_IN;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           TILE2_RXPOLARITY0_IN;
    input           TILE2_RXPOLARITY1_IN;
    //------------------- Shared Ports - Tile and PLL Ports --------------------
    input           TILE2_CLKIN_IN;
    input           TILE2_GTXRESET_IN;
    output          TILE2_PLLLKDET_OUT;
    output          TILE2_REFCLKOUT_OUT;
    output          TILE2_RESETDONE0_OUT;
    output          TILE2_RESETDONE1_OUT;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [19:0]  TILE2_TXDATA0_IN;
    input   [19:0]  TILE2_TXDATA1_IN;
    input           TILE2_TXUSRCLK0_IN;
    input           TILE2_TXUSRCLK1_IN;
    input           TILE2_TXUSRCLK20_IN;
    input           TILE2_TXUSRCLK21_IN;
    //------------- Transmit Ports - TX Driver and OOB signalling --------------
    output          TILE2_TXN0_OUT;
    output          TILE2_TXN1_OUT;
    output          TILE2_TXP0_OUT;
    output          TILE2_TXP1_OUT;





//***************************** Wire Declarations *****************************

    // Channel Bonding Signals




    // ground and vcc signals
    wire            tied_to_ground_i;
    wire    [63:0]  tied_to_ground_vec_i;
    wire            tied_to_vcc_i;
    wire    [63:0]  tied_to_vcc_vec_i;
    
//********************************* Main Body of Code**************************

    assign tied_to_ground_i             = 1'b0;
    assign tied_to_ground_vec_i         = 64'h0000000000000000;
    assign tied_to_vcc_i                = 1'b1;
    assign tied_to_vcc_vec_i            = 64'hffffffffffffffff;
    

    //------------------------- Tile Instances  -------------------------------   



    //_________________________________________________________________________
    //_________________________________________________________________________
    //TILE0  (Location)

    GTX_TILE #
    (
        // Simulation attributes
        .TILE_SIM_MODE               (WRAPPER_SIM_MODE),
        .TILE_SIM_GTXRESET_SPEEDUP   (WRAPPER_SIM_GTXRESET_SPEEDUP),
        .TILE_SIM_PLL_PERDIV2        (WRAPPER_SIM_PLL_PERDIV2),

        // Channel bonding attributes
        .TILE_CHAN_BOND_MODE_0       ("OFF"),
        .TILE_CHAN_BOND_LEVEL_0      (0),
    
        .TILE_CHAN_BOND_MODE_1       ("OFF"),
        .TILE_CHAN_BOND_LEVEL_1      (0)          
    )
    tile0_gtx_i
    (
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
        .RXCHARISCOMMA0_OUT             (TILE0_RXCHARISCOMMA0_OUT),
        .RXCHARISCOMMA1_OUT             (TILE0_RXCHARISCOMMA1_OUT),
        .RXDISPERR0_OUT                 (TILE0_RXDISPERR0_OUT),
        .RXDISPERR1_OUT                 (TILE0_RXDISPERR1_OUT),
        .RXNOTINTABLE0_OUT              (TILE0_RXNOTINTABLE0_OUT),
        .RXNOTINTABLE1_OUT              (TILE0_RXNOTINTABLE1_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXBYTEISALIGNED0_OUT           (TILE0_RXBYTEISALIGNED0_OUT),
        .RXBYTEISALIGNED1_OUT           (TILE0_RXBYTEISALIGNED1_OUT),
        .RXENMCOMMAALIGN0_IN            (TILE0_RXENMCOMMAALIGN0_IN),
        .RXENMCOMMAALIGN1_IN            (TILE0_RXENMCOMMAALIGN1_IN),
        .RXENPCOMMAALIGN0_IN            (TILE0_RXENPCOMMAALIGN0_IN),
        .RXENPCOMMAALIGN1_IN            (TILE0_RXENPCOMMAALIGN1_IN),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .RXDATA0_OUT                    (TILE0_RXDATA0_OUT),
        .RXDATA1_OUT                    (TILE0_RXDATA1_OUT),
        .RXRECCLK0_OUT                  (TILE0_RXRECCLK0_OUT),
        .RXRECCLK1_OUT                  (TILE0_RXRECCLK1_OUT),
        .RXUSRCLK0_IN                   (TILE0_RXUSRCLK0_IN),
        .RXUSRCLK1_IN                   (TILE0_RXUSRCLK1_IN),
        .RXUSRCLK20_IN                  (TILE0_RXUSRCLK20_IN),
        .RXUSRCLK21_IN                  (TILE0_RXUSRCLK21_IN),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .RXEQMIX0_IN                    (TILE0_RXEQMIX0_IN),
        .RXEQMIX1_IN                    (TILE0_RXEQMIX1_IN),
        .RXN0_IN                        (TILE0_RXN0_IN),
        .RXN1_IN                        (TILE0_RXN1_IN),
        .RXP0_IN                        (TILE0_RXP0_IN),
        .RXP1_IN                        (TILE0_RXP1_IN),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY0_IN                 (TILE0_RXPOLARITY0_IN),
        .RXPOLARITY1_IN                 (TILE0_RXPOLARITY1_IN),
        //------------------- Shared Ports - Tile and PLL Ports --------------------
        .CLKIN_IN                       (TILE0_CLKIN_IN),
        .GTXRESET_IN                    (TILE0_GTXRESET_IN),
        .PLLLKDET_OUT                   (TILE0_PLLLKDET_OUT),
        .REFCLKOUT_OUT                  (TILE0_REFCLKOUT_OUT),
        .RESETDONE0_OUT                 (TILE0_RESETDONE0_OUT),
        .RESETDONE1_OUT                 (TILE0_RESETDONE1_OUT),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .TXDATA0_IN                     (TILE0_TXDATA0_IN),
        .TXDATA1_IN                     (TILE0_TXDATA1_IN),
        .TXUSRCLK0_IN                   (TILE0_TXUSRCLK0_IN),
        .TXUSRCLK1_IN                   (TILE0_TXUSRCLK1_IN),
        .TXUSRCLK20_IN                  (TILE0_TXUSRCLK20_IN),
        .TXUSRCLK21_IN                  (TILE0_TXUSRCLK21_IN),
        //------------- Transmit Ports - TX Driver and OOB signalling --------------
        .TXN0_OUT                       (TILE0_TXN0_OUT),
        .TXN1_OUT                       (TILE0_TXN1_OUT),
        .TXP0_OUT                       (TILE0_TXP0_OUT),
        .TXP1_OUT                       (TILE0_TXP1_OUT)

    );



    //_________________________________________________________________________
    //_________________________________________________________________________
    //TILE1  (Location)

    GTX_TILE #
    (
        // Simulation attributes
        .TILE_SIM_MODE               (WRAPPER_SIM_MODE),
        .TILE_SIM_GTXRESET_SPEEDUP   (WRAPPER_SIM_GTXRESET_SPEEDUP),
        .TILE_SIM_PLL_PERDIV2        (WRAPPER_SIM_PLL_PERDIV2),

        // Channel bonding attributes
        .TILE_CHAN_BOND_MODE_0       ("OFF"),
        .TILE_CHAN_BOND_LEVEL_0      (0),
    
        .TILE_CHAN_BOND_MODE_1       ("OFF"),
        .TILE_CHAN_BOND_LEVEL_1      (0)          
    )
    tile1_gtx_i
    (
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
        .RXCHARISCOMMA0_OUT             (TILE1_RXCHARISCOMMA0_OUT),
        .RXCHARISCOMMA1_OUT             (TILE1_RXCHARISCOMMA1_OUT),
        .RXDISPERR0_OUT                 (TILE1_RXDISPERR0_OUT),
        .RXDISPERR1_OUT                 (TILE1_RXDISPERR1_OUT),
        .RXNOTINTABLE0_OUT              (TILE1_RXNOTINTABLE0_OUT),
        .RXNOTINTABLE1_OUT              (TILE1_RXNOTINTABLE1_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXBYTEISALIGNED0_OUT           (TILE1_RXBYTEISALIGNED0_OUT),
        .RXBYTEISALIGNED1_OUT           (TILE1_RXBYTEISALIGNED1_OUT),
        .RXENMCOMMAALIGN0_IN            (TILE1_RXENMCOMMAALIGN0_IN),
        .RXENMCOMMAALIGN1_IN            (TILE1_RXENMCOMMAALIGN1_IN),
        .RXENPCOMMAALIGN0_IN            (TILE1_RXENPCOMMAALIGN0_IN),
        .RXENPCOMMAALIGN1_IN            (TILE1_RXENPCOMMAALIGN1_IN),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .RXDATA0_OUT                    (TILE1_RXDATA0_OUT),
        .RXDATA1_OUT                    (TILE1_RXDATA1_OUT),
        .RXRECCLK0_OUT                  (TILE1_RXRECCLK0_OUT),
        .RXRECCLK1_OUT                  (TILE1_RXRECCLK1_OUT),
        .RXUSRCLK0_IN                   (TILE1_RXUSRCLK0_IN),
        .RXUSRCLK1_IN                   (TILE1_RXUSRCLK1_IN),
        .RXUSRCLK20_IN                  (TILE1_RXUSRCLK20_IN),
        .RXUSRCLK21_IN                  (TILE1_RXUSRCLK21_IN),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .RXEQMIX0_IN                    (TILE1_RXEQMIX0_IN),
        .RXEQMIX1_IN                    (TILE1_RXEQMIX1_IN),
        .RXN0_IN                        (TILE1_RXN0_IN),
        .RXN1_IN                        (TILE1_RXN1_IN),
        .RXP0_IN                        (TILE1_RXP0_IN),
        .RXP1_IN                        (TILE1_RXP1_IN),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY0_IN                 (TILE1_RXPOLARITY0_IN),
        .RXPOLARITY1_IN                 (TILE1_RXPOLARITY1_IN),
        //------------------- Shared Ports - Tile and PLL Ports --------------------
        .CLKIN_IN                       (TILE1_CLKIN_IN),
        .GTXRESET_IN                    (TILE1_GTXRESET_IN),
        .PLLLKDET_OUT                   (TILE1_PLLLKDET_OUT),
        .REFCLKOUT_OUT                  (TILE1_REFCLKOUT_OUT),
        .RESETDONE0_OUT                 (TILE1_RESETDONE0_OUT),
        .RESETDONE1_OUT                 (TILE1_RESETDONE1_OUT),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .TXDATA0_IN                     (TILE1_TXDATA0_IN),
        .TXDATA1_IN                     (TILE1_TXDATA1_IN),
        .TXUSRCLK0_IN                   (TILE1_TXUSRCLK0_IN),
        .TXUSRCLK1_IN                   (TILE1_TXUSRCLK1_IN),
        .TXUSRCLK20_IN                  (TILE1_TXUSRCLK20_IN),
        .TXUSRCLK21_IN                  (TILE1_TXUSRCLK21_IN),
        //------------- Transmit Ports - TX Driver and OOB signalling --------------
        .TXN0_OUT                       (TILE1_TXN0_OUT),
        .TXN1_OUT                       (TILE1_TXN1_OUT),
        .TXP0_OUT                       (TILE1_TXP0_OUT),
        .TXP1_OUT                       (TILE1_TXP1_OUT)

    );



    //_________________________________________________________________________
    //_________________________________________________________________________
    //TILE2  (Location)

    GTX_TILE #
    (
        // Simulation attributes
        .TILE_SIM_MODE               (WRAPPER_SIM_MODE),
        .TILE_SIM_GTXRESET_SPEEDUP   (WRAPPER_SIM_GTXRESET_SPEEDUP),
        .TILE_SIM_PLL_PERDIV2        (WRAPPER_SIM_PLL_PERDIV2),

        // Channel bonding attributes
        .TILE_CHAN_BOND_MODE_0       ("OFF"),
        .TILE_CHAN_BOND_LEVEL_0      (0),
    
        .TILE_CHAN_BOND_MODE_1       ("OFF"),
        .TILE_CHAN_BOND_LEVEL_1      (0)          
    )
    tile2_gtx_i
    (
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
        .RXCHARISCOMMA0_OUT             (TILE2_RXCHARISCOMMA0_OUT),
        .RXCHARISCOMMA1_OUT             (TILE2_RXCHARISCOMMA1_OUT),
        .RXDISPERR0_OUT                 (TILE2_RXDISPERR0_OUT),
        .RXDISPERR1_OUT                 (TILE2_RXDISPERR1_OUT),
        .RXNOTINTABLE0_OUT              (TILE2_RXNOTINTABLE0_OUT),
        .RXNOTINTABLE1_OUT              (TILE2_RXNOTINTABLE1_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXBYTEISALIGNED0_OUT           (TILE2_RXBYTEISALIGNED0_OUT),
        .RXBYTEISALIGNED1_OUT           (TILE2_RXBYTEISALIGNED1_OUT),
        .RXENMCOMMAALIGN0_IN            (TILE2_RXENMCOMMAALIGN0_IN),
        .RXENMCOMMAALIGN1_IN            (TILE2_RXENMCOMMAALIGN1_IN),
        .RXENPCOMMAALIGN0_IN            (TILE2_RXENPCOMMAALIGN0_IN),
        .RXENPCOMMAALIGN1_IN            (TILE2_RXENPCOMMAALIGN1_IN),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .RXDATA0_OUT                    (TILE2_RXDATA0_OUT),
        .RXDATA1_OUT                    (TILE2_RXDATA1_OUT),
        .RXRECCLK0_OUT                  (TILE2_RXRECCLK0_OUT),
        .RXRECCLK1_OUT                  (TILE2_RXRECCLK1_OUT),
        .RXUSRCLK0_IN                   (TILE2_RXUSRCLK0_IN),
        .RXUSRCLK1_IN                   (TILE2_RXUSRCLK1_IN),
        .RXUSRCLK20_IN                  (TILE2_RXUSRCLK20_IN),
        .RXUSRCLK21_IN                  (TILE2_RXUSRCLK21_IN),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .RXEQMIX0_IN                    (TILE2_RXEQMIX0_IN),
        .RXEQMIX1_IN                    (TILE2_RXEQMIX1_IN),
        .RXN0_IN                        (TILE2_RXN0_IN),
        .RXN1_IN                        (TILE2_RXN1_IN),
        .RXP0_IN                        (TILE2_RXP0_IN),
        .RXP1_IN                        (TILE2_RXP1_IN),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY0_IN                 (TILE2_RXPOLARITY0_IN),
        .RXPOLARITY1_IN                 (TILE2_RXPOLARITY1_IN),
        //------------------- Shared Ports - Tile and PLL Ports --------------------
        .CLKIN_IN                       (TILE2_CLKIN_IN),
        .GTXRESET_IN                    (TILE2_GTXRESET_IN),
        .PLLLKDET_OUT                   (TILE2_PLLLKDET_OUT),
        .REFCLKOUT_OUT                  (TILE2_REFCLKOUT_OUT),
        .RESETDONE0_OUT                 (TILE2_RESETDONE0_OUT),
        .RESETDONE1_OUT                 (TILE2_RESETDONE1_OUT),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .TXDATA0_IN                     (TILE2_TXDATA0_IN),
        .TXDATA1_IN                     (TILE2_TXDATA1_IN),
        .TXUSRCLK0_IN                   (TILE2_TXUSRCLK0_IN),
        .TXUSRCLK1_IN                   (TILE2_TXUSRCLK1_IN),
        .TXUSRCLK20_IN                  (TILE2_TXUSRCLK20_IN),
        .TXUSRCLK21_IN                  (TILE2_TXUSRCLK21_IN),
        //------------- Transmit Ports - TX Driver and OOB signalling --------------
        .TXN0_OUT                       (TILE2_TXN0_OUT),
        .TXN1_OUT                       (TILE2_TXN1_OUT),
        .TXP0_OUT                       (TILE2_TXP0_OUT),
        .TXP1_OUT                       (TILE2_TXP1_OUT)

    );

    
     
endmodule

