///////////////////////////////////////////////////////////////////////////////
//$Date: 2008/07/23 00:15:51 $
//$RCSfile: example_mgt_top.ejava,v $
//$Revision: 1.1.2.6 $
////////////////////////////////////////////////////////////////////////////////
//   ____  ____ 
//  /   /\/   / 
// /___/  \  /    Vendor: Xilinx 
// \   \   \/     Version : 1.5
//  \   \         Application : GTX Wizard 
//  /   /         Filename : example_mgt_top.v
// /___/   /\     Timestamp : 
// \   \  /  \ 
//  \___\/\___\ 
//
//
// Module EXAMPLE_MGT_TOP
// Generated by Xilinx GTX Wizard




`timescale 1ns / 1ps
`define DLY #1


//***********************************Entity Declaration************************

module EXAMPLE_MGT_TOP #
(
    parameter EXAMPLE_CONFIG_INDEPENDENT_LANES          =   1,   //configuration for frame gen and check
    parameter EXAMPLE_LANE_WITH_START_CHAR              =   0,   // specifies lane with unique start frame char
    parameter EXAMPLE_WORDS_IN_BRAM                     =   512, // specifies amount of data in BRAM 
    parameter EXAMPLE_SIM_MODE                          =   "FAST",  // Set to Fast Functional Simulation Model
    parameter EXAMPLE_SIM_GTXRESET_SPEEDUP              =   1,   // simulation setting for MGT smartmodel
    parameter EXAMPLE_SIM_PLL_PERDIV2                   =   9'h0fa, // simulation setting for MGT smartmodel
    parameter EXAMPLE_USE_CHIPSCOPE                     =   1    // Set to 1 to use Chipscope to drive resets
)
(
    GREFCLK_N_IN,
    GREFCLK_P_IN,
    GTXRESET_IN,
    TILE0_PLLLKDET_OUT,
    TILE1_PLLLKDET_OUT,
    RXN_IN,
    RXP_IN,
    TXN_OUT,
    TXP_OUT
);

// synthesis attribute X_CORE_INFO of EXAMPLE_MGT_TOP is "gtxwizard_v1_5, Coregen v10.1_ip3";

//***********************************Ports Declaration*******************************

    input           GREFCLK_N_IN;
    input           GREFCLK_P_IN;
    input           GTXRESET_IN;
    output          TILE0_PLLLKDET_OUT;
    output          TILE1_PLLLKDET_OUT;
    input   [3:0]   RXN_IN;
    input   [3:0]   RXP_IN;
    output  [3:0]   TXN_OUT;
    output  [3:0]   TXP_OUT;

    
//************************** Register Declarations ****************************

    reg     [84:0]  ila_in0_r;
    reg     [84:0]  ila_in1_r;
    reg             tile0_tx_resetdone0_r;
    reg             tile0_tx_resetdone0_r2;
    reg             tile0_rx_resetdone0_r;
    reg             tile0_rx_resetdone0_r2;
    reg             tile0_tx_resetdone1_r;
    reg             tile0_tx_resetdone1_r2;
    reg             tile0_rx_resetdone1_r;
    reg             tile0_rx_resetdone1_r2;
    reg             tile1_tx_resetdone0_r;
    reg             tile1_tx_resetdone0_r2;
    reg             tile1_rx_resetdone0_r;
    reg             tile1_rx_resetdone0_r2;
    reg             tile1_tx_resetdone1_r;
    reg             tile1_tx_resetdone1_r2;
    reg             tile1_rx_resetdone1_r;
    reg             tile1_rx_resetdone1_r2;
    

//**************************** Wire Declarations ******************************

    //------------------------ MGT Wrapper Wires ------------------------------
    

    //________________________________________________________________________
    //________________________________________________________________________
    //TILE0   (X0Y3)

    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    wire    [1:0]   tile0_rxchariscomma0_i;
    wire    [1:0]   tile0_rxchariscomma1_i;
    wire    [1:0]   tile0_rxdisperr0_i;
    wire    [1:0]   tile0_rxdisperr1_i;
    wire    [1:0]   tile0_rxnotintable0_i;
    wire    [1:0]   tile0_rxnotintable1_i;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    wire            tile0_rxbyteisaligned0_i;
    wire            tile0_rxbyteisaligned1_i;
    wire            tile0_rxbyterealign0_i;
    wire            tile0_rxbyterealign1_i;
    wire            tile0_rxenmcommaalign0_i;
    wire            tile0_rxenmcommaalign1_i;
    wire            tile0_rxenpcommaalign0_i;
    wire            tile0_rxenpcommaalign1_i;
    //----------------- Receive Ports - RX Data Path interface -----------------
    wire    [15:0]  tile0_rxdata0_i;
    wire    [15:0]  tile0_rxdata1_i;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    wire    [1:0]   tile0_rxeqmix0_i;
    wire    [1:0]   tile0_rxeqmix1_i;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    wire            tile0_rxpolarity0_i;
    wire            tile0_rxpolarity1_i;
    //------------------- Shared Ports - Tile and PLL Ports --------------------
    wire            tile0_gtxreset_i;
    wire            tile0_plllkdet_i;
    wire            tile0_refclkout_i;
    wire            tile0_resetdone0_i;
    wire            tile0_resetdone1_i;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    wire    [19:0]  tile0_txdata0_i;
    wire    [19:0]  tile0_txdata1_i;



    //________________________________________________________________________
    //________________________________________________________________________
    //TILE1   (X0Y5)

    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    wire    [1:0]   tile1_rxchariscomma0_i;
    wire    [1:0]   tile1_rxchariscomma1_i;
    wire    [1:0]   tile1_rxdisperr0_i;
    wire    [1:0]   tile1_rxdisperr1_i;
    wire    [1:0]   tile1_rxnotintable0_i;
    wire    [1:0]   tile1_rxnotintable1_i;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    wire            tile1_rxbyteisaligned0_i;
    wire            tile1_rxbyteisaligned1_i;
    wire            tile1_rxbyterealign0_i;
    wire            tile1_rxbyterealign1_i;
    wire            tile1_rxenmcommaalign0_i;
    wire            tile1_rxenmcommaalign1_i;
    wire            tile1_rxenpcommaalign0_i;
    wire            tile1_rxenpcommaalign1_i;
    //----------------- Receive Ports - RX Data Path interface -----------------
    wire    [15:0]  tile1_rxdata0_i;
    wire    [15:0]  tile1_rxdata1_i;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    wire    [1:0]   tile1_rxeqmix0_i;
    wire    [1:0]   tile1_rxeqmix1_i;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    wire            tile1_rxpolarity0_i;
    wire            tile1_rxpolarity1_i;
    //------------------- Shared Ports - Tile and PLL Ports --------------------
    wire            tile1_gtxreset_i;
    wire            tile1_plllkdet_i;
    wire            tile1_refclkout_i;
    wire            tile1_resetdone0_i;
    wire            tile1_resetdone1_i;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    wire    [19:0]  tile1_txdata0_i;
    wire    [19:0]  tile1_txdata1_i;


    //----------------------------- Global Signals -----------------------------
    wire            tile0_tx_system_reset0_c;
    wire            tile0_rx_system_reset0_c;
    wire            tile0_tx_system_reset1_c;
    wire            tile0_rx_system_reset1_c;
    wire            tile1_tx_system_reset0_c;
    wire            tile1_rx_system_reset0_c;
    wire            tile1_tx_system_reset1_c;
    wire            tile1_rx_system_reset1_c;
    wire            tied_to_ground_i;
    wire    [63:0]  tied_to_ground_vec_i;
    wire            tied_to_vcc_i;
    wire    [7:0]   tied_to_vcc_vec_i;
    wire            drp_clk_in_i;
    wire            grefclk_i;
    
    wire            tile0_refclkout_bufg_i;
    
    
    //--------------------------- User Clocks ---------------------------------
    wire            tile0_txusrclk0_i;


    //--------------------- Frame check/gen Module Signals --------------------
    wire            tile0_matchn0_i;
    
    wire    [1:0]   tile0_txcharisk0_float_i;
    
    wire    [19:0]  tile0_txdata0_float_i;
    
    
    wire            tile0_block_sync0_reset_i;
    wire    [7:0]   tile0_error_count0_i;
    wire            tile0_frame_check0_reset_i;
    wire            tile0_inc_in0_i;
    wire            tile0_inc_out0_i;
    wire    [15:0]  tile0_unscrambled_data0_i;
    wire            tile0_matchn1_i;
    
    wire    [1:0]   tile0_txcharisk1_float_i;
    
    wire    [19:0]  tile0_txdata1_float_i;
    
    
    wire            tile0_block_sync1_reset_i;
    wire    [7:0]   tile0_error_count1_i;
    wire            tile0_frame_check1_reset_i;
    wire            tile0_inc_in1_i;
    wire            tile0_inc_out1_i;
    wire    [15:0]  tile0_unscrambled_data1_i;

    wire            tile1_matchn0_i;
    
    wire    [1:0]   tile1_txcharisk0_float_i;
    
    wire    [19:0]  tile1_txdata0_float_i;
    
    
    wire            tile1_block_sync0_reset_i;
    wire    [7:0]   tile1_error_count0_i;
    wire            tile1_frame_check0_reset_i;
    wire            tile1_inc_in0_i;
    wire            tile1_inc_out0_i;
    wire    [15:0]  tile1_unscrambled_data0_i;
    wire            tile1_matchn1_i;
    
    wire    [1:0]   tile1_txcharisk1_float_i;
    
    wire    [19:0]  tile1_txdata1_float_i;
    
    
    wire            tile1_block_sync1_reset_i;
    wire    [7:0]   tile1_error_count1_i;
    wire            tile1_frame_check1_reset_i;
    wire            tile1_inc_in1_i;
    wire            tile1_inc_out1_i;
    wire    [15:0]  tile1_unscrambled_data1_i;

    wire            reset_on_data_error_i;
    wire            grefclk_in_i;


    //--------------------- Chipscope Signals ---------------------------------

    wire    [35:0]  shared_vio_control_i;
    wire    [35:0]  tx_data_vio_control0_i;
    wire    [35:0]  tx_data_vio_control1_i;
    wire    [35:0]  rx_data_vio_control0_i;
    wire    [35:0]  rx_data_vio_control1_i;
    wire    [35:0]  ila_control0_i;
    wire    [35:0]  ila_control1_i;
    wire    [31:0]  shared_vio_in_i;
    wire    [31:0]  shared_vio_out_i;
    wire    [31:0]  tx_data_vio_in0_i;
    wire    [31:0]  tx_data_vio_out0_i;
    wire    [31:0]  tx_data_vio_in1_i;
    wire    [31:0]  tx_data_vio_out1_i;
    wire    [31:0]  rx_data_vio_in0_i;
    wire    [31:0]  rx_data_vio_out0_i;
    wire    [31:0]  rx_data_vio_in1_i;
    wire    [31:0]  rx_data_vio_out1_i;
    wire    [84:0]  ila_in0_i;
    wire    [84:0]  ila_in1_i;

    wire    [31:0]  tile0_tx_data_vio_in0_i;
    wire    [31:0]  tile0_tx_data_vio_out0_i;
    wire    [31:0]  tile0_tx_data_vio_in1_i;
    wire    [31:0]  tile0_tx_data_vio_out1_i;
    wire    [31:0]  tile0_rx_data_vio_in0_i;
    wire    [31:0]  tile0_rx_data_vio_out0_i;
    wire    [31:0]  tile0_rx_data_vio_in1_i;
    wire    [31:0]  tile0_rx_data_vio_out1_i;
    wire    [84:0]  tile0_ila_in0_i;
    wire    [84:0]  tile0_ila_in1_i;

    wire    [31:0]  tile1_tx_data_vio_in0_i;
    wire    [31:0]  tile1_tx_data_vio_out0_i;
    wire    [31:0]  tile1_tx_data_vio_in1_i;
    wire    [31:0]  tile1_tx_data_vio_out1_i;
    wire    [31:0]  tile1_rx_data_vio_in0_i;
    wire    [31:0]  tile1_rx_data_vio_out0_i;
    wire    [31:0]  tile1_rx_data_vio_in1_i;
    wire    [31:0]  tile1_rx_data_vio_out1_i;
    wire    [84:0]  tile1_ila_in0_i;
    wire    [84:0]  tile1_ila_in1_i;


    wire            gtxreset_i;
    wire            mux_sel_i;
    wire            user_tx_reset_i;
    wire            user_rx_reset_i;
    wire            ila_clk0_i;
    wire            ila_clk_mux_out0_i;
    wire            ila_clk1_i;
    wire            ila_clk_mux_out1_i;


//**************************** Main Body of Code *******************************

    //  Static signal Assigments    
    assign tied_to_ground_i             = 1'b0;
    assign tied_to_ground_vec_i         = 64'h0000000000000000;
    assign tied_to_vcc_i                = 1'b1;
    assign tied_to_vcc_vec_i            = 8'hff;


    






    //----- Reference clock using normal clock resources (GREFCLK)  -----------
    // In designs that can tolerate higher jitter, GREFCLK reference clock inputs to the GTXs can
    // be used. In this example, we use an IBUFDS to bring a reference clock on chip through the
    // regular IOs    
        
    IBUFDS grefclk_ibufds_i
    (
        .O                              (grefclk_in_i), 
        .I                              (GREFCLK_P_IN),
        .IB                             (GREFCLK_N_IN)
    );

    // The tools automatically turn on GREFCLK reference clocking when the CLKIN port of the GTX is 
    // driven by a BUFG. Here we connect the grefclk from the IBUFDS to a BUFG, which we will use to 
    // drive the GTXs in the design that were selected to use GREFCLK.
    
    BUFG grefclk_bufg_i
    (
        .I                              (grefclk_in_i),
        .O                              (grefclk_i) 
    );



    //--------------------------------- User Clocks ---------------------------
    
    // The clock resources in this section were added based on userclk source selections on
    // the Latency, Buffering, and Clocking page of the GUI. A few notes about user clocks:
    // * The userclk and userclk2 for each GTX datapath (TX and RX) must be phase aligned to 
    //   avoid data errors in the fabric interface whenever the datapath is wider than 10 bits
    // * To minimize clock resources, you can share clocks between GTXs. GTXs using the same frequency
    //   or multiples of the same frequency can be accomadated using DCMs and PLLs. Use caution when
    //   using RXRECCLK as a clock source, however - these clocks can typically only be shared if all
    //   the channels using the clock are receiving data from TX channels that share a reference clock 
    //   source with each other.

    BUFG refclkout_bufg0_i
    (
        .I                              (tile0_refclkout_i),
        .O                              (tile0_txusrclk0_i)
    );






    //--------------------------- The GTX Wrapper -----------------------------
    
    // Use the instantiation template in the examples directory to add the GTX wrapper to your design.
    // In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    // checker. The GTXs will reset, then attempt to align and transmit data. If channel bonding is 
    // enabled, bonding should occur after alignment.
 
    
    // Wire all PLLLKDET signals to the top level as output ports
    assign TILE0_PLLLKDET_OUT = tile0_plllkdet_i;
    assign TILE1_PLLLKDET_OUT = tile1_plllkdet_i;


    GTX #
    (
        .WRAPPER_SIM_MODE               (EXAMPLE_SIM_MODE),
        .WRAPPER_SIM_GTXRESET_SPEEDUP   (EXAMPLE_SIM_GTXRESET_SPEEDUP),
        .WRAPPER_SIM_PLL_PERDIV2        (EXAMPLE_SIM_PLL_PERDIV2)
    )
    gtx_i
    (
    
 
 
 
 
 
 
 
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //TILE0  (X0Y3)

        //--------------------- Receive Ports - 8b10b Decoder ----------------------
        .TILE0_RXCHARISCOMMA0_OUT       (tile0_rxchariscomma0_i),
        .TILE0_RXCHARISCOMMA1_OUT       (tile0_rxchariscomma1_i),
        .TILE0_RXDISPERR0_OUT           (tile0_rxdisperr0_i),
        .TILE0_RXDISPERR1_OUT           (tile0_rxdisperr1_i),
        .TILE0_RXNOTINTABLE0_OUT        (tile0_rxnotintable0_i),
        .TILE0_RXNOTINTABLE1_OUT        (tile0_rxnotintable1_i),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .TILE0_RXBYTEISALIGNED0_OUT     (tile0_rxbyteisaligned0_i),
        .TILE0_RXBYTEISALIGNED1_OUT     (tile0_rxbyteisaligned1_i),
        .TILE0_RXBYTEREALIGN0_OUT       (tile0_rxbyterealign0_i),
        .TILE0_RXBYTEREALIGN1_OUT       (tile0_rxbyterealign1_i),
        .TILE0_RXENMCOMMAALIGN0_IN      (tile0_rxenmcommaalign0_i),
        .TILE0_RXENMCOMMAALIGN1_IN      (tile0_rxenmcommaalign1_i),
        .TILE0_RXENPCOMMAALIGN0_IN      (tile0_rxenpcommaalign0_i),
        .TILE0_RXENPCOMMAALIGN1_IN      (tile0_rxenpcommaalign1_i),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .TILE0_RXDATA0_OUT              (tile0_rxdata0_i),
        .TILE0_RXDATA1_OUT              (tile0_rxdata1_i),
        .TILE0_RXUSRCLK0_IN             (tile0_txusrclk0_i),
        .TILE0_RXUSRCLK1_IN             (tile0_txusrclk0_i),
        .TILE0_RXUSRCLK20_IN            (tile0_txusrclk0_i),
        .TILE0_RXUSRCLK21_IN            (tile0_txusrclk0_i),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .TILE0_RXEQMIX0_IN              (tile0_rxeqmix0_i),
        .TILE0_RXEQMIX1_IN              (tile0_rxeqmix1_i),
        .TILE0_RXN0_IN                  (RXN_IN[0]),
        .TILE0_RXN1_IN                  (RXN_IN[1]),
        .TILE0_RXP0_IN                  (RXP_IN[0]),
        .TILE0_RXP1_IN                  (RXP_IN[1]),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .TILE0_RXPOLARITY0_IN           (tile0_rxpolarity0_i),
        .TILE0_RXPOLARITY1_IN           (tile0_rxpolarity1_i),
        //------------------- Shared Ports - Tile and PLL Ports --------------------
        .TILE0_CLKIN_IN                 (grefclk_i),
        .TILE0_GTXRESET_IN              (tile0_gtxreset_i),
        .TILE0_PLLLKDET_OUT             (tile0_plllkdet_i),
        .TILE0_REFCLKOUT_OUT            (tile0_refclkout_i),
        .TILE0_RESETDONE0_OUT           (tile0_resetdone0_i),
        .TILE0_RESETDONE1_OUT           (tile0_resetdone1_i),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .TILE0_TXDATA0_IN               (tile0_txdata0_i),
        .TILE0_TXDATA1_IN               (tile0_txdata1_i),
        .TILE0_TXUSRCLK0_IN             (tile0_txusrclk0_i),
        .TILE0_TXUSRCLK1_IN             (tile0_txusrclk0_i),
        .TILE0_TXUSRCLK20_IN            (tile0_txusrclk0_i),
        .TILE0_TXUSRCLK21_IN            (tile0_txusrclk0_i),
        //------------- Transmit Ports - TX Driver and OOB signalling --------------
        .TILE0_TXN0_OUT                 (TXN_OUT[0]),
        .TILE0_TXN1_OUT                 (TXN_OUT[1]),
        .TILE0_TXP0_OUT                 (TXP_OUT[0]),
        .TILE0_TXP1_OUT                 (TXP_OUT[1]),


    
 
 
 
 
 
 
 
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //TILE1  (X0Y5)

        //--------------------- Receive Ports - 8b10b Decoder ----------------------
        .TILE1_RXCHARISCOMMA0_OUT       (tile1_rxchariscomma0_i),
        .TILE1_RXCHARISCOMMA1_OUT       (tile1_rxchariscomma1_i),
        .TILE1_RXDISPERR0_OUT           (tile1_rxdisperr0_i),
        .TILE1_RXDISPERR1_OUT           (tile1_rxdisperr1_i),
        .TILE1_RXNOTINTABLE0_OUT        (tile1_rxnotintable0_i),
        .TILE1_RXNOTINTABLE1_OUT        (tile1_rxnotintable1_i),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .TILE1_RXBYTEISALIGNED0_OUT     (tile1_rxbyteisaligned0_i),
        .TILE1_RXBYTEISALIGNED1_OUT     (tile1_rxbyteisaligned1_i),
        .TILE1_RXBYTEREALIGN0_OUT       (tile1_rxbyterealign0_i),
        .TILE1_RXBYTEREALIGN1_OUT       (tile1_rxbyterealign1_i),
        .TILE1_RXENMCOMMAALIGN0_IN      (tile1_rxenmcommaalign0_i),
        .TILE1_RXENMCOMMAALIGN1_IN      (tile1_rxenmcommaalign1_i),
        .TILE1_RXENPCOMMAALIGN0_IN      (tile1_rxenpcommaalign0_i),
        .TILE1_RXENPCOMMAALIGN1_IN      (tile1_rxenpcommaalign1_i),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .TILE1_RXDATA0_OUT              (tile1_rxdata0_i),
        .TILE1_RXDATA1_OUT              (tile1_rxdata1_i),
        .TILE1_RXUSRCLK0_IN             (tile0_txusrclk0_i),
        .TILE1_RXUSRCLK1_IN             (tile0_txusrclk0_i),
        .TILE1_RXUSRCLK20_IN            (tile0_txusrclk0_i),
        .TILE1_RXUSRCLK21_IN            (tile0_txusrclk0_i),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .TILE1_RXEQMIX0_IN              (tile1_rxeqmix0_i),
        .TILE1_RXEQMIX1_IN              (tile1_rxeqmix1_i),
        .TILE1_RXN0_IN                  (RXN_IN[2]),
        .TILE1_RXN1_IN                  (RXN_IN[3]),
        .TILE1_RXP0_IN                  (RXP_IN[2]),
        .TILE1_RXP1_IN                  (RXP_IN[3]),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .TILE1_RXPOLARITY0_IN           (tile1_rxpolarity0_i),
        .TILE1_RXPOLARITY1_IN           (tile1_rxpolarity1_i),
        //------------------- Shared Ports - Tile and PLL Ports --------------------
        .TILE1_CLKIN_IN                 (grefclk_i),
        .TILE1_GTXRESET_IN              (tile1_gtxreset_i),
        .TILE1_PLLLKDET_OUT             (tile1_plllkdet_i),
        .TILE1_REFCLKOUT_OUT            (tile1_refclkout_i),
        .TILE1_RESETDONE0_OUT           (tile1_resetdone0_i),
        .TILE1_RESETDONE1_OUT           (tile1_resetdone1_i),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .TILE1_TXDATA0_IN               (tile1_txdata0_i),
        .TILE1_TXDATA1_IN               (tile1_txdata1_i),
        .TILE1_TXUSRCLK0_IN             (tile0_txusrclk0_i),
        .TILE1_TXUSRCLK1_IN             (tile0_txusrclk0_i),
        .TILE1_TXUSRCLK20_IN            (tile0_txusrclk0_i),
        .TILE1_TXUSRCLK21_IN            (tile0_txusrclk0_i),
        //------------- Transmit Ports - TX Driver and OOB signalling --------------
        .TILE1_TXN0_OUT                 (TXN_OUT[2]),
        .TILE1_TXN1_OUT                 (TXN_OUT[3]),
        .TILE1_TXP0_OUT                 (TXP_OUT[2]),
        .TILE1_TXP1_OUT                 (TXP_OUT[3])


    );







    //------------------------ User Module Resets -----------------------------
    // All the User Modules i.e. FRAME_GEN, FRAME_CHECK and the sync modules
    // are held in reset till the RESETDONE goes high. 
    // The RESETDONE is registered a couple of times on *USRCLK2 and connected 
    // to the reset of the modules
    
    always @(posedge tile0_txusrclk0_i or negedge tile0_resetdone0_i)

    begin
        if (!tile0_resetdone0_i )
        begin
            tile0_rx_resetdone0_r    <=   `DLY 1'b0;
            tile0_rx_resetdone0_r2   <=   `DLY 1'b0;
        end
        else
        begin
            tile0_rx_resetdone0_r    <=   `DLY tile0_resetdone0_i;
            tile0_rx_resetdone0_r2   <=   `DLY tile0_rx_resetdone0_r;
        end
    end
    
    
    always @(posedge tile0_txusrclk0_i or negedge tile0_resetdone0_i)

    begin
        if (!tile0_resetdone0_i )
        begin
            tile0_tx_resetdone0_r    <=   `DLY 1'b0;
            tile0_tx_resetdone0_r2   <=   `DLY 1'b0;
        end
        else
        begin
            tile0_tx_resetdone0_r    <=   `DLY tile0_resetdone0_i;
            tile0_tx_resetdone0_r2   <=   `DLY tile0_tx_resetdone0_r;
        end
    end
    always @(posedge tile0_txusrclk0_i or negedge tile0_resetdone1_i)

    begin
        if (!tile0_resetdone1_i )
        begin
            tile0_rx_resetdone1_r    <=   `DLY 1'b0;
            tile0_rx_resetdone1_r2   <=   `DLY 1'b0;
        end
        else
        begin
            tile0_rx_resetdone1_r    <=   `DLY tile0_resetdone1_i;
            tile0_rx_resetdone1_r2   <=   `DLY tile0_rx_resetdone1_r;
        end
    end
    
    
    always @(posedge tile0_txusrclk0_i or negedge tile0_resetdone1_i)

    begin
        if (!tile0_resetdone1_i )
        begin
            tile0_tx_resetdone1_r    <=   `DLY 1'b0;
            tile0_tx_resetdone1_r2   <=   `DLY 1'b0;
        end
        else
        begin
            tile0_tx_resetdone1_r    <=   `DLY tile0_resetdone1_i;
            tile0_tx_resetdone1_r2   <=   `DLY tile0_tx_resetdone1_r;
        end
    end
    always @(posedge tile0_txusrclk0_i or negedge tile1_resetdone0_i)

    begin
        if (!tile1_resetdone0_i )
        begin
            tile1_rx_resetdone0_r    <=   `DLY 1'b0;
            tile1_rx_resetdone0_r2   <=   `DLY 1'b0;
        end
        else
        begin
            tile1_rx_resetdone0_r    <=   `DLY tile1_resetdone0_i;
            tile1_rx_resetdone0_r2   <=   `DLY tile1_rx_resetdone0_r;
        end
    end
    
    
    always @(posedge tile0_txusrclk0_i or negedge tile1_resetdone0_i)

    begin
        if (!tile1_resetdone0_i )
        begin
            tile1_tx_resetdone0_r    <=   `DLY 1'b0;
            tile1_tx_resetdone0_r2   <=   `DLY 1'b0;
        end
        else
        begin
            tile1_tx_resetdone0_r    <=   `DLY tile1_resetdone0_i;
            tile1_tx_resetdone0_r2   <=   `DLY tile1_tx_resetdone0_r;
        end
    end
    always @(posedge tile0_txusrclk0_i or negedge tile1_resetdone1_i)

    begin
        if (!tile1_resetdone1_i )
        begin
            tile1_rx_resetdone1_r    <=   `DLY 1'b0;
            tile1_rx_resetdone1_r2   <=   `DLY 1'b0;
        end
        else
        begin
            tile1_rx_resetdone1_r    <=   `DLY tile1_resetdone1_i;
            tile1_rx_resetdone1_r2   <=   `DLY tile1_rx_resetdone1_r;
        end
    end
    
    
    always @(posedge tile0_txusrclk0_i or negedge tile1_resetdone1_i)

    begin
        if (!tile1_resetdone1_i )
        begin
            tile1_tx_resetdone1_r    <=   `DLY 1'b0;
            tile1_tx_resetdone1_r2   <=   `DLY 1'b0;
        end
        else
        begin
            tile1_tx_resetdone1_r    <=   `DLY tile1_resetdone1_i;
            tile1_tx_resetdone1_r2   <=   `DLY tile1_tx_resetdone1_r;
        end
    end

    



    //---------------------------- Frame Generators ---------------------------
    // The example design uses Block RAM based frame generators to provide test
    // data to the GTXs for transmission. By default the frame generators are 
    // loaded with an incrementing data sequence that includes commas/alignment
    // characters for alignment. If your protocol uses channel bonding, the 
    // frame generator will also be preloaded with a channel bonding sequence.
    
    // You can modify the data transmitted by changing the INIT values of the frame
    // generator in this file. Pay careful attention to bit order and the spacing
    // of your control and alignment characters.

    FRAME_GEN #
    (
        .WORDS_IN_BRAM(EXAMPLE_WORDS_IN_BRAM),
        .MEM_00(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_01(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_02(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_03(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_04(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_05(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_06(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_07(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_08(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_09(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_0A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_0B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_0C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_0D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_0E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_0F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_10(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_11(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_12(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_13(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_14(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_15(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_16(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_17(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_18(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_19(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_1A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_1B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_1C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_1D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_1E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_1F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_20(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_21(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_22(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_23(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_24(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_25(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_26(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_27(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_28(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_29(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_2A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_2B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_2C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_2D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_2E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_2F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_30(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_31(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_32(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_33(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_34(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_35(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_36(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_37(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_38(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_39(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_3A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_3B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_3C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_3D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_3E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_3F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEMP_00(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_01(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_02(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_03(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_04(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_05(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_06(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_07(256'h0000000000000000000000000000000000000000000000000000000000000010)
    )
    tile0_frame_gen0
    (
        // User Interface
        .TX_DATA                        ({tile0_txdata0_float_i,tile0_txdata0_i}),
    
        .TX_CHARISK                     ( ),
        // System Interface
        .USER_CLK                       (tile0_txusrclk0_i),
        .SYSTEM_RESET                   (tile0_tx_system_reset0_c)
    );

    FRAME_GEN #
    (
        .WORDS_IN_BRAM(EXAMPLE_WORDS_IN_BRAM),
        .MEM_00(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_01(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_02(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_03(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_04(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_05(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_06(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_07(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_08(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_09(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_0A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_0B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_0C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_0D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_0E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_0F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_10(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_11(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_12(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_13(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_14(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_15(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_16(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_17(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_18(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_19(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_1A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_1B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_1C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_1D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_1E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_1F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_20(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_21(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_22(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_23(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_24(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_25(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_26(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_27(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_28(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_29(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_2A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_2B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_2C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_2D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_2E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_2F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_30(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_31(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_32(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_33(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_34(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_35(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_36(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_37(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_38(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_39(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_3A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_3B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_3C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_3D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_3E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_3F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEMP_00(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_01(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_02(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_03(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_04(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_05(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_06(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_07(256'h0000000000000000000000000000000000000000000000000000000000000010)
    )
    tile0_frame_gen1
    (
        // User Interface
        .TX_DATA                        ({tile0_txdata1_float_i,tile0_txdata1_i}),
    
        .TX_CHARISK                     ( ),
        // System Interface
        .USER_CLK                       (tile0_txusrclk0_i),
        .SYSTEM_RESET                   (tile0_tx_system_reset1_c)
    );

    FRAME_GEN #
    (
        .WORDS_IN_BRAM(EXAMPLE_WORDS_IN_BRAM),
        .MEM_00(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_01(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_02(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_03(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_04(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_05(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_06(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_07(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_08(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_09(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_0A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_0B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_0C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_0D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_0E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_0F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_10(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_11(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_12(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_13(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_14(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_15(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_16(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_17(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_18(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_19(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_1A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_1B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_1C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_1D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_1E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_1F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_20(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_21(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_22(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_23(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_24(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_25(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_26(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_27(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_28(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_29(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_2A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_2B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_2C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_2D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_2E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_2F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_30(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_31(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_32(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_33(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_34(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_35(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_36(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_37(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_38(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_39(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_3A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_3B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_3C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_3D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_3E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_3F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEMP_00(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_01(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_02(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_03(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_04(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_05(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_06(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_07(256'h0000000000000000000000000000000000000000000000000000000000000010)
    )
    tile1_frame_gen0
    (
        // User Interface
        .TX_DATA                        ({tile1_txdata0_float_i,tile1_txdata0_i}),
    
        .TX_CHARISK                     ( ),
        // System Interface
        .USER_CLK                       (tile0_txusrclk0_i),
        .SYSTEM_RESET                   (tile1_tx_system_reset0_c)
    );

    FRAME_GEN #
    (
        .WORDS_IN_BRAM(EXAMPLE_WORDS_IN_BRAM),
        .MEM_00(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_01(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_02(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_03(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_04(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_05(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_06(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_07(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_08(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_09(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_0A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_0B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_0C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_0D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_0E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_0F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_10(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_11(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_12(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_13(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_14(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_15(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_16(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_17(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_18(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_19(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_1A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_1B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_1C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_1D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_1E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_1F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_20(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_21(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_22(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_23(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_24(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_25(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_26(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_27(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_28(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_29(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_2A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_2B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_2C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_2D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_2E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_2F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_30(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_31(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_32(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_33(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_34(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_35(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_36(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_37(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEM_38(256'h0000380d0000300b00002809000020070000180500001003000002bc00000400),
        .MEM_39(256'h0000781d0000701b00006819000060170000581500005013000048110000400f),
        .MEM_3A(256'h0000b82d0000b02b0000a8290000a0270000982500009023000088210000801f),
        .MEM_3B(256'h0000f83d0000f03b0000e8390000e0370000d8350000d0330000c8310000c02f),
        .MEM_3C(256'h0001384d0001304b00012849000120470001184500011043000108410001003f),
        .MEM_3D(256'h0001785d0001705b00016859000160570001585500015053000148510001404f),
        .MEM_3E(256'h0001b86d0001b06b0001a8690001a0670001986500019063000188610001805f),
        .MEM_3F(256'h0001f87d0001f07b0001e8790001e0770001d8750001d0730001c8710001c06f),
        .MEMP_00(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_01(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_02(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_03(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_04(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_05(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_06(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_07(256'h0000000000000000000000000000000000000000000000000000000000000010)
    )
    tile1_frame_gen1
    (
        // User Interface
        .TX_DATA                        ({tile1_txdata1_float_i,tile1_txdata1_i}),
    
        .TX_CHARISK                     ( ),
        // System Interface
        .USER_CLK                       (tile0_txusrclk0_i),
        .SYSTEM_RESET                   (tile1_tx_system_reset1_c)
    );



    //-------------------------------- Frame Checkers -------------------------
    // The example design uses Block RAM based frame checkers to verify incoming  
    // data. By default the frame generators are loaded with a data sequence that 
    // matches the outgoing sequence of the frame generators for the TX ports.
    
    // You can modify the expected data sequence by changing the INIT values of the frame
    // checkers in this file. Pay careful attention to bit order and the spacing
    // of your control and alignment characters.
    
    // When the frame checker receives data, it attempts to synchronise to the 
    // incoming pattern by looking for the first sequence in the pattern. Once it 
    // finds the first sequence, it increments through the sequence, and indicates an 
    // error whenever the next value received does not match the expected value.


    assign tile0_frame_check0_reset_i = (EXAMPLE_CONFIG_INDEPENDENT_LANES==0)?reset_on_data_error_i:tile0_matchn0_i;

    // tile0_frame_check0 is always connected to the lane with the start of char
    // and this lane starts off the data checking on all the other lanes. The INC_IN port is tied off
    assign tile0_inc_in0_i = 1'b0;

    FRAME_CHECK #
    (
        .RX_DATA_WIDTH(16),
        .USE_COMMA(1),
        .WORDS_IN_BRAM(EXAMPLE_WORDS_IN_BRAM),
        .CONFIG_INDEPENDENT_LANES(1),
        .START_OF_PACKET_CHAR(8'hbc),
        .MEM_00(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_01(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_02(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_03(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_04(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_05(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_06(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_07(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_08(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_09(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_0A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_0B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_0C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_0D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_0E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_0F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_10(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_11(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_12(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_13(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_14(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_15(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_16(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_17(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_18(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_19(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_1A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_1B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_1C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_1D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_1E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_1F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_20(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_21(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_22(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_23(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_24(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_25(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_26(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_27(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_28(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_29(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_2A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_2B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_2C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_2D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_2E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_2F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_30(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_31(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_32(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_33(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_34(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_35(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_36(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_37(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_38(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_39(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_3A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_3B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_3C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_3D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_3E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_3F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEMP_00(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_01(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_02(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_03(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_04(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_05(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_06(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_07(256'h0000000000000000000000000000000000000000000000000000000000000010)
    )
    tile0_frame_check0
    (
        // MGT Interface
        .RX_DATA                        (tile0_rxdata0_i),  
        .RX_ENMCOMMA_ALIGN              (tile0_rxenmcommaalign0_i),
        .RX_ENPCOMMA_ALIGN              (tile0_rxenpcommaalign0_i),
        .RX_ENCHAN_SYNC                 ( ),
        .RX_CHANBOND_SEQ                (tied_to_ground_i),
        // Control Interface
        .INC_IN                         (tile0_inc_in0_i),
        .INC_OUT                        (tile0_inc_out0_i),
        .PATTERN_MATCH_N                (tile0_matchn0_i),
        .RESET_ON_ERROR                 (tile0_frame_check0_reset_i),
        // System Interface
        .USER_CLK                       (tile0_txusrclk0_i),
        .SYSTEM_RESET                   (tile0_rx_system_reset0_c),
        .ERROR_COUNT                    (tile0_error_count0_i)
  
    );

    

    assign tile0_frame_check1_reset_i = (EXAMPLE_CONFIG_INDEPENDENT_LANES==0)?reset_on_data_error_i:tile0_matchn1_i;

    // tile0_frame_check0 is always connected to the lane with the start of char
    // and this lane starts off the data checking on all the other lanes. The INC_IN port is tied off
    assign tile0_inc_in1_i = 1'b0;

    FRAME_CHECK #
    (
        .RX_DATA_WIDTH(16),
        .USE_COMMA(1),
        .WORDS_IN_BRAM(EXAMPLE_WORDS_IN_BRAM),
        .CONFIG_INDEPENDENT_LANES(1),
        .START_OF_PACKET_CHAR(8'hbc),
        .MEM_00(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_01(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_02(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_03(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_04(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_05(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_06(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_07(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_08(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_09(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_0A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_0B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_0C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_0D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_0E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_0F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_10(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_11(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_12(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_13(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_14(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_15(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_16(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_17(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_18(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_19(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_1A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_1B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_1C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_1D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_1E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_1F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_20(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_21(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_22(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_23(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_24(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_25(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_26(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_27(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_28(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_29(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_2A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_2B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_2C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_2D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_2E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_2F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_30(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_31(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_32(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_33(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_34(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_35(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_36(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_37(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_38(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_39(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_3A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_3B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_3C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_3D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_3E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_3F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEMP_00(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_01(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_02(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_03(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_04(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_05(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_06(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_07(256'h0000000000000000000000000000000000000000000000000000000000000010)
    )
    tile0_frame_check1
    (
        // MGT Interface
        .RX_DATA                        (tile0_rxdata1_i),  
        .RX_ENMCOMMA_ALIGN              (tile0_rxenmcommaalign1_i),
        .RX_ENPCOMMA_ALIGN              (tile0_rxenpcommaalign1_i),
        .RX_ENCHAN_SYNC                 ( ),
        .RX_CHANBOND_SEQ                (tied_to_ground_i),
        // Control Interface
        .INC_IN                         (tile0_inc_in1_i),
        .INC_OUT                        (tile0_inc_out1_i),
        .PATTERN_MATCH_N                (tile0_matchn1_i),
        .RESET_ON_ERROR                 (tile0_frame_check1_reset_i),
        // System Interface
        .USER_CLK                       (tile0_txusrclk0_i),
        .SYSTEM_RESET                   (tile0_rx_system_reset1_c),
        .ERROR_COUNT                    (tile0_error_count1_i)
  
    );

    

    assign tile1_frame_check0_reset_i = (EXAMPLE_CONFIG_INDEPENDENT_LANES==0)?reset_on_data_error_i:tile1_matchn0_i;

    // in the "independent lanes" configuration, each of the lanes looks for the unique start char and
    // in this case, the INC_IN port is tied off.
    // Else, the data checking is triggered by the "master" lane
    assign tile1_inc_in0_i = (EXAMPLE_CONFIG_INDEPENDENT_LANES==0)?tile0_inc_out0_i:1'b0;

    FRAME_CHECK #
    (
        .RX_DATA_WIDTH(16),
        .USE_COMMA(1),
        .WORDS_IN_BRAM(EXAMPLE_WORDS_IN_BRAM),
        .CONFIG_INDEPENDENT_LANES(EXAMPLE_CONFIG_INDEPENDENT_LANES),
        .START_OF_PACKET_CHAR(8'hbc),
        .MEM_00(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_01(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_02(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_03(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_04(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_05(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_06(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_07(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_08(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_09(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_0A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_0B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_0C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_0D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_0E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_0F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_10(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_11(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_12(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_13(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_14(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_15(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_16(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_17(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_18(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_19(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_1A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_1B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_1C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_1D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_1E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_1F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_20(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_21(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_22(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_23(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_24(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_25(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_26(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_27(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_28(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_29(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_2A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_2B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_2C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_2D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_2E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_2F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_30(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_31(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_32(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_33(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_34(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_35(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_36(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_37(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_38(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_39(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_3A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_3B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_3C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_3D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_3E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_3F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEMP_00(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_01(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_02(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_03(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_04(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_05(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_06(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_07(256'h0000000000000000000000000000000000000000000000000000000000000010)
    )
    tile1_frame_check0
    (
        // MGT Interface
        .RX_DATA                        (tile1_rxdata0_i),  
        .RX_ENMCOMMA_ALIGN              (tile1_rxenmcommaalign0_i),
        .RX_ENPCOMMA_ALIGN              (tile1_rxenpcommaalign0_i),
        .RX_ENCHAN_SYNC                 ( ),
        .RX_CHANBOND_SEQ                (tied_to_ground_i),
        // Control Interface
        .INC_IN                         (tile1_inc_in0_i),
        .INC_OUT                        (tile1_inc_out0_i),
        .PATTERN_MATCH_N                (tile1_matchn0_i),
        .RESET_ON_ERROR                 (tile1_frame_check0_reset_i),
        // System Interface
        .USER_CLK                       (tile0_txusrclk0_i),
        .SYSTEM_RESET                   (tile1_rx_system_reset0_c),
        .ERROR_COUNT                    (tile1_error_count0_i)
  
    );

    

    assign tile1_frame_check1_reset_i = (EXAMPLE_CONFIG_INDEPENDENT_LANES==0)?reset_on_data_error_i:tile1_matchn1_i;

    // in the "independent lanes" configuration, each of the lanes looks for the unique start char and
    // in this case, the INC_IN port is tied off.
    // Else, the data checking is triggered by the "master" lane
    assign tile1_inc_in1_i = (EXAMPLE_CONFIG_INDEPENDENT_LANES==0)?tile0_inc_out1_i:1'b0;

    FRAME_CHECK #
    (
        .RX_DATA_WIDTH(16),
        .USE_COMMA(1),
        .WORDS_IN_BRAM(EXAMPLE_WORDS_IN_BRAM),
        .CONFIG_INDEPENDENT_LANES(EXAMPLE_CONFIG_INDEPENDENT_LANES),
        .START_OF_PACKET_CHAR(8'hbc),
        .MEM_00(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_01(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_02(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_03(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_04(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_05(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_06(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_07(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_08(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_09(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_0A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_0B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_0C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_0D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_0E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_0F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_10(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_11(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_12(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_13(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_14(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_15(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_16(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_17(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_18(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_19(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_1A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_1B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_1C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_1D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_1E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_1F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_20(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_21(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_22(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_23(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_24(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_25(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_26(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_27(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_28(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_29(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_2A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_2B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_2C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_2D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_2E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_2F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_30(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_31(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_32(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_33(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_34(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_35(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_36(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_37(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEM_38(256'h00000e0d00000c0b00000a09000008070000060500000403000002bc00000100),
        .MEM_39(256'h00001e1d00001c1b00001a19000018170000161500001413000012110000100f),
        .MEM_3A(256'h00002e2d00002c2b00002a29000028270000262500002423000022210000201f),
        .MEM_3B(256'h00003e3d00003c3b00003a39000038370000363500003433000032310000302f),
        .MEM_3C(256'h00004e4d00004c4b00004a49000048470000464500004443000042410000403f),
        .MEM_3D(256'h00005e5d00005c5b00005a59000058570000565500005453000052510000504f),
        .MEM_3E(256'h00006e6d00006c6b00006a69000068670000666500006463000062610000605f),
        .MEM_3F(256'h00007e7d00007c7b00007a79000078770000767500007473000072710000706f),
        .MEMP_00(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_01(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_02(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_03(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_04(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_05(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_06(256'h0000000000000000000000000000000000000000000000000000000000000010),
        .MEMP_07(256'h0000000000000000000000000000000000000000000000000000000000000010)
    )
    tile1_frame_check1
    (
        // MGT Interface
        .RX_DATA                        (tile1_rxdata1_i),  
        .RX_ENMCOMMA_ALIGN              (tile1_rxenmcommaalign1_i),
        .RX_ENPCOMMA_ALIGN              (tile1_rxenpcommaalign1_i),
        .RX_ENCHAN_SYNC                 ( ),
        .RX_CHANBOND_SEQ                (tied_to_ground_i),
        // Control Interface
        .INC_IN                         (tile1_inc_in1_i),
        .INC_OUT                        (tile1_inc_out1_i),
        .PATTERN_MATCH_N                (tile1_matchn1_i),
        .RESET_ON_ERROR                 (tile1_frame_check1_reset_i),
        // System Interface
        .USER_CLK                       (tile0_txusrclk0_i),
        .SYSTEM_RESET                   (tile1_rx_system_reset1_c),
        .ERROR_COUNT                    (tile1_error_count1_i)
  
    );

    





    //--------------------------- Chipscope Connections -----------------------
    // When the example design is run in hardware, it uses chipscope to allow the
    // example design and GTX wrapper to be controlled and monitored. The 
    // EXAMPLE_USE_CHIPSCOPE parameter allows chipscope to be removed for simulation.
    
generate
if (EXAMPLE_USE_CHIPSCOPE==1) 
begin : chipscope


    // Shared VIO for all tiles
    shared_vio shared_vio_i
    (
      .control                          (shared_vio_control_i),
      .async_in                         (shared_vio_in_i),
      .async_out                        (shared_vio_out_i)
    );

    // ICON for all VIOs 
    icon i_icon
    (
      .control0                         (shared_vio_control_i),
      .control1                         (tx_data_vio_control0_i),
      .control2                         (rx_data_vio_control0_i),
      .control3                         (ila_control0_i),
      .control4                         (tx_data_vio_control1_i),
      .control5                         (rx_data_vio_control1_i),
      .control6                         (ila_control1_i)
    );

    // TX VIO 
    shared_vio tx_data_vio0_i
    (
      .control                          (tx_data_vio_control0_i),
      .async_in                         (tx_data_vio_in0_i),
      .async_out                        (tx_data_vio_out0_i)  
    );
    
    // RX VIO 
    shared_vio rx_data_vio0_i
    (
      .control                          (rx_data_vio_control0_i),
      .async_in                         (rx_data_vio_in0_i),
      .async_out                        (rx_data_vio_out0_i)  
    );
    
    // RX ILA
    ila ila0_i
    (
      .control                          (ila_control0_i),
      .clk                              (ila_clk0_i),
      .trig0                            (ila_in0_i)
    );


    
    // The RX ILA must use the same clock as the selected transceiver
    BUFG ila_clk0_bufg_i
    (
        .I      (ila_clk_mux_out0_i),
        .O      (ila_clk0_i)
    );

    assign  ila_clk_mux_out0_i = tile0_txusrclk0_i;


    // TX VIO 
    shared_vio tx_data_vio1_i
    (
      .control                          (tx_data_vio_control1_i),
      .async_in                         (tx_data_vio_in1_i),
      .async_out                        (tx_data_vio_out1_i)  
    );
    
    // RX VIO 
    shared_vio rx_data_vio1_i
    (
      .control                          (rx_data_vio_control1_i),
      .async_in                         (rx_data_vio_in1_i),
      .async_out                        (rx_data_vio_out1_i)  
    );
    
    // RX ILA
    ila ila1_i
    (
      .control                          (ila_control1_i),
      .clk                              (ila_clk1_i),
      .trig0                            (ila_in1_i)
    );


    
    // The RX ILA must use the same clock as the selected transceiver
    BUFG ila_clk1_bufg_i
    (
        .I      (ila_clk_mux_out1_i),
        .O      (ila_clk1_i)
    );

    assign  ila_clk_mux_out1_i = tile0_txusrclk0_i;



    // assign resets for frame_gen modules
    assign  tile0_tx_system_reset0_c = !tile0_tx_resetdone0_r2 || user_tx_reset_i;
    assign  tile0_tx_system_reset1_c = !tile0_tx_resetdone1_r2 || user_tx_reset_i;
    assign  tile1_tx_system_reset0_c = !tile1_tx_resetdone0_r2 || user_tx_reset_i;
    assign  tile1_tx_system_reset1_c = !tile1_tx_resetdone1_r2 || user_tx_reset_i;

    // assign resets for frame_check modules
    assign  tile0_rx_system_reset0_c = !tile0_rx_resetdone0_r2 || user_rx_reset_i;
    assign  tile0_rx_system_reset1_c = !tile0_rx_resetdone1_r2 || user_rx_reset_i;
    assign  tile1_rx_system_reset0_c = !tile1_rx_resetdone0_r2 || user_rx_reset_i;
    assign  tile1_rx_system_reset1_c = !tile1_rx_resetdone1_r2 || user_rx_reset_i;


    assign  tile0_gtxreset_i = gtxreset_i;
    assign  tile1_gtxreset_i = gtxreset_i;

    // Shared VIO Outputs
    assign  gtxreset_i                      =  shared_vio_out_i[31];
    assign  user_tx_reset_i                 =  shared_vio_out_i[30];
    assign  user_rx_reset_i                 =  shared_vio_out_i[29];
    assign  mux_sel_i                       =  shared_vio_out_i[28];

    // Shared VIO Inputs
    assign  shared_vio_in_i[31]             =  tile0_plllkdet_i;
    assign  shared_vio_in_i[30]             =  tile1_plllkdet_i;
    assign  shared_vio_in_i[29:0]           =  30'b000000000000000000000000000000;

    // Chipscope connections for GTP0 on Tile 0
    assign  tile0_tx_data_vio_in0_i[31:0]   =  32'b00000000000000000000000000000000;
    assign  tile0_rx_data_vio_in0_i[31]     =  tile0_resetdone0_i;
    assign  tile0_rx_data_vio_in0_i[30:0]   =  31'b0000000000000000000000000000000;
    assign  tile0_rxeqmix0_i                =  rx_data_vio_out0_i[31:30];
    assign  tile0_rxpolarity0_i             =  rx_data_vio_out0_i[29];
    assign  tile0_ila_in0_i[84:83]          =  tile0_rxchariscomma0_i;
    assign  tile0_ila_in0_i[82:81]          =  tile0_rxdisperr0_i;
    assign  tile0_ila_in0_i[80:79]          =  tile0_rxnotintable0_i;
    assign  tile0_ila_in0_i[78]             =  tile0_rxbyteisaligned0_i;
    assign  tile0_ila_in0_i[77]             =  tile0_rxbyterealign0_i;
    assign  tile0_ila_in0_i[76:61]          =  tile0_rxdata0_i;
    assign  tile0_ila_in0_i[60:53]          =  tile0_error_count0_i;
    assign  tile0_ila_in0_i[52:0]           =  53'b00000000000000000000000000000000000000000000000000000;

    // Chipscope connections for GTP1 on Tile 0
    assign  tile0_tx_data_vio_in1_i[31:0]   =  32'b00000000000000000000000000000000;
    assign  tile0_rx_data_vio_in1_i[31]     =  tile0_resetdone1_i;
    assign  tile0_rx_data_vio_in1_i[30:0]   =  31'b0000000000000000000000000000000;
    assign  tile0_rxeqmix1_i                =  rx_data_vio_out1_i[31:30];
    assign  tile0_rxpolarity1_i             =  rx_data_vio_out1_i[29];
    assign  tile0_ila_in1_i[84:83]          =  tile0_rxchariscomma1_i;
    assign  tile0_ila_in1_i[82:81]          =  tile0_rxdisperr1_i;
    assign  tile0_ila_in1_i[80:79]          =  tile0_rxnotintable1_i;
    assign  tile0_ila_in1_i[78]             =  tile0_rxbyteisaligned1_i;
    assign  tile0_ila_in1_i[77]             =  tile0_rxbyterealign1_i;
    assign  tile0_ila_in1_i[76:61]          =  tile0_rxdata1_i;
    assign  tile0_ila_in1_i[60:53]          =  tile0_error_count1_i;
    assign  tile0_ila_in1_i[52:0]           =  53'b00000000000000000000000000000000000000000000000000000;

    // Chipscope connections for GTP0 on Tile 1
    assign  tile1_tx_data_vio_in0_i[31:0]   =  32'b00000000000000000000000000000000;
    assign  tile1_rx_data_vio_in0_i[31]     =  tile1_resetdone0_i;
    assign  tile1_rx_data_vio_in0_i[30:0]   =  31'b0000000000000000000000000000000;
    assign  tile1_rxeqmix0_i                =  rx_data_vio_out0_i[31:30];
    assign  tile1_rxpolarity0_i             =  rx_data_vio_out0_i[29];
    assign  tile1_ila_in0_i[84:83]          =  tile1_rxchariscomma0_i;
    assign  tile1_ila_in0_i[82:81]          =  tile1_rxdisperr0_i;
    assign  tile1_ila_in0_i[80:79]          =  tile1_rxnotintable0_i;
    assign  tile1_ila_in0_i[78]             =  tile1_rxbyteisaligned0_i;
    assign  tile1_ila_in0_i[77]             =  tile1_rxbyterealign0_i;
    assign  tile1_ila_in0_i[76:61]          =  tile1_rxdata0_i;
    assign  tile1_ila_in0_i[60:53]          =  tile1_error_count0_i;
    assign  tile1_ila_in0_i[52:0]           =  53'b00000000000000000000000000000000000000000000000000000;

    // Chipscope connections for GTP1 on Tile 1
    assign  tile1_tx_data_vio_in1_i[31:0]   =  32'b00000000000000000000000000000000;
    assign  tile1_rx_data_vio_in1_i[31]     =  tile1_resetdone1_i;
    assign  tile1_rx_data_vio_in1_i[30:0]   =  31'b0000000000000000000000000000000;
    assign  tile1_rxeqmix1_i                =  rx_data_vio_out1_i[31:30];
    assign  tile1_rxpolarity1_i             =  rx_data_vio_out1_i[29];
    assign  tile1_ila_in1_i[84:83]          =  tile1_rxchariscomma1_i;
    assign  tile1_ila_in1_i[82:81]          =  tile1_rxdisperr1_i;
    assign  tile1_ila_in1_i[80:79]          =  tile1_rxnotintable1_i;
    assign  tile1_ila_in1_i[78]             =  tile1_rxbyteisaligned1_i;
    assign  tile1_ila_in1_i[77]             =  tile1_rxbyterealign1_i;
    assign  tile1_ila_in1_i[76:61]          =  tile1_rxdata1_i;
    assign  tile1_ila_in1_i[60:53]          =  tile1_error_count1_i;
    assign  tile1_ila_in1_i[52:0]           =  53'b00000000000000000000000000000000000000000000000000000;


    //Mux inputs to Chipscope modules based on mux_sel_i

    assign  tx_data_vio_in0_i =         (mux_sel_i == 1'b0)?tile0_tx_data_vio_in0_i:
                                                            tile1_tx_data_vio_in0_i;


    assign  rx_data_vio_in0_i =         (mux_sel_i == 1'b0)?tile0_rx_data_vio_in0_i:
                                                            tile1_rx_data_vio_in0_i;


    assign  ila_in0_i =                 (mux_sel_i == 1'b0)?tile0_ila_in0_i:
                                                            tile1_ila_in0_i;


    assign  tx_data_vio_in1_i =         (mux_sel_i == 1'b0)?tile0_tx_data_vio_in1_i:
                                                            tile1_tx_data_vio_in1_i;


    assign  rx_data_vio_in1_i =         (mux_sel_i == 1'b0)?tile0_rx_data_vio_in1_i:
                                                            tile1_rx_data_vio_in1_i;


    assign  ila_in1_i =                 (mux_sel_i == 1'b0)?tile0_ila_in1_i:
                                                            tile1_ila_in1_i;




end //end EXAMPLE_USE_CHIPSCOPE=1 generate section
else 
begin: no_chipscope

    // If Chipscope is not being used, drive GTX reset signal
    // from the top level ports
    assign  tile0_gtxreset_i = GTXRESET_IN;
    assign  tile1_gtxreset_i = GTXRESET_IN;

    // assign resets for frame_gen modules
    assign  tile0_tx_system_reset0_c = !tile0_tx_resetdone0_r2;
    assign  tile0_tx_system_reset1_c = !tile0_tx_resetdone1_r2;
    assign  tile1_tx_system_reset0_c = !tile1_tx_resetdone0_r2;
    assign  tile1_tx_system_reset1_c = !tile1_tx_resetdone1_r2;

    // assign resets for frame_check modules
    assign  tile0_rx_system_reset0_c = !tile0_rx_resetdone0_r2;
    assign  tile0_rx_system_reset1_c = !tile0_rx_resetdone1_r2;
    assign  tile1_rx_system_reset0_c = !tile1_rx_resetdone0_r2;
    assign  tile1_rx_system_reset1_c = !tile1_rx_resetdone1_r2;

    assign  gtxreset_i                      =  tied_to_ground_i;
    assign  user_tx_reset_i                 =  tied_to_ground_i;
    assign  user_rx_reset_i                 =  tied_to_ground_i;
    assign  mux_sel_i                       =  tied_to_ground_i;
    assign  tile0_rxeqmix0_i                =  tied_to_ground_vec_i[1:0];
    assign  tile0_rxpolarity0_i             =  tied_to_ground_i;
    assign  tile0_rxeqmix1_i                =  tied_to_ground_vec_i[1:0];
    assign  tile0_rxpolarity1_i             =  tied_to_ground_i;
    assign  tile1_rxeqmix0_i                =  tied_to_ground_vec_i[1:0];
    assign  tile1_rxpolarity0_i             =  tied_to_ground_i;
    assign  tile1_rxeqmix1_i                =  tied_to_ground_vec_i[1:0];
    assign  tile1_rxpolarity1_i             =  tied_to_ground_i;



end
endgenerate //End generate for EXAMPLE_USE_CHIPSCOPE


endmodule

//-------------------------------------------------------------------
//
//  VIO core module declaration 
//  This one is for driving shared ports and is asynchronous
//
//-------------------------------------------------------------------
module shared_vio
  (
    control,
    async_in,
    async_out
  );
  input  [35:0] control;
  input  [31:0] async_in;
  output [31:0] async_out;
endmodule

//-------------------------------------------------------------------
//
//  ICON core module declaration
//
//-------------------------------------------------------------------
module icon
  (
      control0,
      control1,
      control2,
      control3,
      control4,
      control5,
      control6  );
  output [35:0] control0;
  output [35:0] control1;
  output [35:0] control2;
  output [35:0] control3;
  output [35:0] control4;
  output [35:0] control5;
  output [35:0] control6;
endmodule


//-------------------------------------------------------------------
//
//  ILA core module declaration
//  This is used to allow RX signals to be monitored
//
//-------------------------------------------------------------------
module ila
  (
    control,
    clk,
    trig0
  );
  input [35:0] control;
  input clk;
  input [84:0] trig0;
endmodule


