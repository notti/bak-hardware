-------------------------------------------------------------------------------
--$Date: 2008/05/30 00:57:53 $
--$RCSfile: example_tb_vhd.ejava,v $
--$Revision: 1.1.2.1 $
--------------------------------------------------------------------------------
--   ____  ____ 
--  /   /\/   / 
-- /___/  \  /    Vendor: Xilinx 
-- \   \   \/     Version : 1.5
--  \   \         Application : RocketIO GTX Wizard 
--  /   /         Filename : example_tb.vhd
-- /___/   /\     Timestamp : 
-- \   \  /  \ 
--  \___\/\___\ 
--
--
-- Module EXAMPLE_TB
-- Generated by Xilinx RocketIO GTX Wizard
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

entity EXAMPLE_TB is
end EXAMPLE_TB;

architecture RTL of EXAMPLE_TB is

--*************************Parameter Declarations******************************

    constant   REFCLK_PERIOD        :   time :=  10.0 ns;
  
--**************************** Component Declarations *************************

    component EXAMPLE_MGT_TOP 
    generic
    (
        EXAMPLE_CONFIG_INDEPENDENT_LANES: integer    := 1;
        EXAMPLE_LANE_WITH_START_CHAR    : integer    := 0;
        EXAMPLE_WORDS_IN_BRAM           : integer    := 512;
        EXAMPLE_SIM_MODE                : string     := "FAST";
        EXAMPLE_SIM_GTXRESET_SPEEDUP    : integer    := 1;
        EXAMPLE_SIM_PLL_PERDIV2         : bit_vector := x"0fa";
        EXAMPLE_USE_CHIPSCOPE           : integer    := 0     --0 - drive resets from top level ports
    );
    port
    (
        TILE2_REFCLK_PAD_N_IN   :   in std_logic;
        TILE2_REFCLK_PAD_P_IN   :   in std_logic; 
        GTXRESET_IN                       :   in std_logic; 
        TILE0_PLLLKDET_OUT                :   out std_logic;
        TILE1_PLLLKDET_OUT                :   out std_logic;
        TILE2_PLLLKDET_OUT                :   out std_logic;
        RXN_IN                            :   in std_logic_vector(5 downto 0);
        RXP_IN                            :   in std_logic_vector(5 downto 0);
        TXN_OUT                           :   out std_logic_vector(5 downto 0);
        TXP_OUT                           :   out std_logic_vector(5 downto 0)
    );
    end component;

    component SIM_RESET_MGT_MODEL 
    port 
    (
        GSR_IN     : in std_logic
    );
    end component;

--************************Internal Register Declarations***********************

--************************** Register Declarations ****************************        

    signal  debounce_pma_reset_r    :   std_logic_vector(0 to 3);
    signal  refclk_n_r              :   std_logic;
    signal  drp_clk_r               :   std_logic;
    signal  tx_usrclk_r             :   std_logic;
    signal  rx_usrclk_r             :   std_logic;    
    signal  gsr_r                   :   std_logic;
    signal  gts_r                   :   std_logic;
    signal  reset_i                 :   std_logic;

--********************************Wire Declarations**********************************
    
    ----------------------------------- Global Signals ------------------------------
    signal  refclk_p_r              :   std_logic;
    signal  tied_to_ground_i        :   std_logic;
    ---------------------------- Example Module Connections -------------------------
    signal  rxn_in_i                :   std_logic_vector(5 downto 0);
    signal  rxp_in_i                :   std_logic_vector(5 downto 0);
    signal  txn_out_i               :   std_logic_vector(5 downto 0);
    signal  txp_out_i               :   std_logic_vector(5 downto 0);


    signal  tile0_error_count0_i   :   std_logic_vector(7 downto 0);
    signal  tile0_error_count1_i   :   std_logic_vector(7 downto 0);
    signal  tile0_plllkdet_i       :   std_logic;
    signal  tile1_error_count0_i   :   std_logic_vector(7 downto 0);
    signal  tile1_error_count1_i   :   std_logic_vector(7 downto 0);
    signal  tile1_plllkdet_i       :   std_logic;
    signal  tile2_error_count0_i   :   std_logic_vector(7 downto 0);
    signal  tile2_error_count1_i   :   std_logic_vector(7 downto 0);
    signal  tile2_plllkdet_i       :   std_logic;

    

--*********************************Main Body of Code**********************************
begin

    -- ------------------------------- Tie offs ------------------------------- 
    
    tied_to_ground_i        <=  '0';
    
    -- ------------------------- MGT Serial Connections -----------------------

    rxn_in_i                <=  txn_out_i;
    rxp_in_i                <=  txp_out_i;  

    ------- Instantiate the ROC module for resetting the VHDL MGT Smart Model ------

    sim_reset_mgt_model_i : SIM_RESET_MGT_MODEL  
    port map    
    (
        GSR_IN           =>           reset_i
    );

    ---------------------- Generate Reference Clock input  --------------------
    
    process
    begin
        refclk_n_r  <=  '1';
        wait for REFCLK_PERIOD/2;
        refclk_n_r  <=  '0';
        wait for REFCLK_PERIOD/2;
    end process;

    refclk_p_r <= not refclk_n_r;
                 

 
                
    ----------------------------------- Resets ---------------------------------
    
    process
    begin
        reset_i <= '1';
        wait for 100 ns;
        reset_i <= '0';
        wait; 
    end process;

    ------------------- Instantiate an EXAMPLE_MGT_TOP module  -----------------

    example_mgt_top_i : EXAMPLE_MGT_TOP
    generic map
    (
        EXAMPLE_SIM_MODE            =>  "FAST",     -- Set to Fast Functional Simulation Model
        EXAMPLE_SIM_GTXRESET_SPEEDUP=>  1,        -- Speedup is turned on for simulation
        EXAMPLE_SIM_PLL_PERDIV2     =>  x"0fa",      -- Set to the VCO Unit Interval time
        EXAMPLE_USE_CHIPSCOPE       =>  0         --1 - use chipscope to drive resets,
                                                          --0 - drive resets from top level ports
    )
    port map
    (
        TILE2_REFCLK_PAD_N_IN       =>  refclk_n_r,   
        TILE2_REFCLK_PAD_P_IN       =>  refclk_p_r,
        GTXRESET_IN                 =>  reset_i,
        TILE0_PLLLKDET_OUT          =>  tile0_plllkdet_i,
        TILE1_PLLLKDET_OUT          =>  tile1_plllkdet_i,
        TILE2_PLLLKDET_OUT          =>  tile2_plllkdet_i,
        RXN_IN                      =>  rxn_in_i,
        RXP_IN                      =>  rxp_in_i,
        TXN_OUT                     =>  txn_out_i,
        TXP_OUT                     =>  txp_out_i
    );


end RTL;

